module module_output_bit_63(i,o);

input [1893:0] i;
output  o;

wire [0:0] l_0;
wire [1:0] l_1;
wire [3:0] l_2;
wire [7:0] l_3;
wire [13:0] l_4;
wire [13:0] l_5;
wire [13:0] l_6;
wire [13:0] l_7;
wire [19:0] l_8;
wire [17:0] l_9;
wire [17:0] l_10;

assign	l_10[17:0]	= 18'b0;

assign o = l_0[0];

assign l_0[0]    = ( l_1 [0] & !i[63]) | ( l_1 [1] &  i[63]);
assign l_1[0]    = ( l_2 [0] & !i[1713]) | ( l_2 [1] &  i[1713]);
assign l_1[1]    = ( l_2 [2] & !i[1713]) | ( l_2 [3] &  i[1713]);
assign l_2[0]    = ( l_3 [0] & !i[1714]) | ( l_3 [1] &  i[1714]);
assign l_2[1]    = ( l_3 [2] & !i[1714]) | ( l_3 [3] &  i[1714]);
assign l_2[2]    = ( l_3 [4] & !i[1714]) | ( l_3 [5] &  i[1714]);
assign l_2[3]    = ( l_3 [6] & !i[1714]) | ( l_3 [7] &  i[1714]);
assign l_3[0]    = ( l_4 [0] &  i[1715]);
assign l_3[1]    = ( l_4 [1] & !i[1715]) | ( l_4 [2] &  i[1715]);
assign l_3[2]    = ( l_4 [3] & !i[1715]) | ( l_4 [4] &  i[1715]);
assign l_3[3]    = ( l_4 [5] & !i[1715]) | ( l_4 [6] &  i[1715]);
assign l_3[4]    = (!i[1715]) | ( l_4 [7] &  i[1715]);
assign l_3[5]    = ( l_4 [8] & !i[1715]) | ( l_4 [9] &  i[1715]);
assign l_3[6]    = ( l_4 [10] & !i[1715]) | ( l_4 [11] &  i[1715]);
assign l_3[7]    = ( l_4 [12] & !i[1715]) | ( l_4 [13] &  i[1715]);
assign l_4[0]    = ( l_5 [0] & !i[1716]);
assign l_4[1]    = ( l_5 [1] & !i[1716]);
assign l_4[2]    = ( l_5 [2] & !i[1716]);
assign l_4[3]    = ( l_5 [3] & !i[1716]);
assign l_4[4]    = ( l_5 [4] & !i[1716]);
assign l_4[5]    = ( l_5 [5] & !i[1716]);
assign l_4[6]    = ( l_5 [6] & !i[1716]);
assign l_4[7]    = ( l_5 [7] & !i[1716]) | (      i[1716]);
assign l_4[8]    = ( l_5 [8] & !i[1716]) | (      i[1716]);
assign l_4[9]    = ( l_5 [9] & !i[1716]) | (      i[1716]);
assign l_4[10]    = ( l_5 [10] & !i[1716]) | (      i[1716]);
assign l_4[11]    = ( l_5 [11] & !i[1716]) | (      i[1716]);
assign l_4[12]    = ( l_5 [12] & !i[1716]) | (      i[1716]);
assign l_4[13]    = ( l_5 [13] & !i[1716]) | (      i[1716]);
assign l_5[0]    = ( l_6 [0] & !i[1717]);
assign l_5[1]    = ( l_6 [1] & !i[1717]);
assign l_5[2]    = ( l_6 [2] & !i[1717]);
assign l_5[3]    = ( l_6 [3] & !i[1717]);
assign l_5[4]    = ( l_6 [4] & !i[1717]);
assign l_5[5]    = ( l_6 [5] & !i[1717]);
assign l_5[6]    = ( l_6 [6] & !i[1717]);
assign l_5[7]    = ( l_6 [7] & !i[1717]) | (      i[1717]);
assign l_5[8]    = ( l_6 [8] & !i[1717]) | (      i[1717]);
assign l_5[9]    = ( l_6 [9] & !i[1717]) | (      i[1717]);
assign l_5[10]    = ( l_6 [10] & !i[1717]) | (      i[1717]);
assign l_5[11]    = ( l_6 [11] & !i[1717]) | (      i[1717]);
assign l_5[12]    = ( l_6 [12] & !i[1717]) | (      i[1717]);
assign l_5[13]    = ( l_6 [13] & !i[1717]) | (      i[1717]);
assign l_6[0]    = ( l_7 [0] &  i[1723]);
assign l_6[1]    = ( l_7 [1] &  i[1723]);
assign l_6[2]    = ( l_7 [2] &  i[1723]);
assign l_6[3]    = ( l_7 [3] &  i[1723]);
assign l_6[4]    = ( l_7 [4] &  i[1723]);
assign l_6[5]    = ( l_7 [5] &  i[1723]);
assign l_6[6]    = ( l_7 [6] &  i[1723]);
assign l_6[7]    = (!i[1723]) | ( l_7 [7] &  i[1723]);
assign l_6[8]    = (!i[1723]) | ( l_7 [8] &  i[1723]);
assign l_6[9]    = (!i[1723]) | ( l_7 [9] &  i[1723]);
assign l_6[10]    = (!i[1723]) | ( l_7 [10] &  i[1723]);
assign l_6[11]    = (!i[1723]) | ( l_7 [11] &  i[1723]);
assign l_6[12]    = (!i[1723]) | ( l_7 [12] &  i[1723]);
assign l_6[13]    = (!i[1723]) | ( l_7 [13] &  i[1723]);
assign l_7[0]    = ( l_8 [0] & !i[1707]);
assign l_7[1]    = ( l_8 [1] & !i[1707]) | ( l_8 [2] &  i[1707]);
assign l_7[2]    = ( l_8 [3] & !i[1707]) | ( l_8 [4] &  i[1707]);
assign l_7[3]    = ( l_8 [5] & !i[1707]) | ( l_8 [6] &  i[1707]);
assign l_7[4]    = ( l_8 [7] & !i[1707]) | ( l_8 [8] &  i[1707]);
assign l_7[5]    = ( l_8 [5] & !i[1707]) | ( l_8 [9] &  i[1707]);
assign l_7[6]    = ( l_8 [5] &  i[1707]);
assign l_7[7]    = ( l_8 [10] & !i[1707]) | ( l_8 [11] &  i[1707]);
assign l_7[8]    = ( l_8 [12] & !i[1707]) | ( l_8 [13] &  i[1707]);
assign l_7[9]    = ( l_8 [14] & !i[1707]) | ( l_8 [15] &  i[1707]);
assign l_7[10]    = (!l_8 [6] & !i[1707]) | ( l_8 [16] &  i[1707]);
assign l_7[11]    = ( l_8 [17] & !i[1707]) | ( l_8 [18] &  i[1707]);
assign l_7[12]    = (!l_8 [6] & !i[1707]) | (      i[1707]);
assign l_7[13]    = (!l_8 [9] & !i[1707]) | ( l_8 [19] &  i[1707]);
assign l_8[0]    = ( l_9 [0] & !i[1724]);
assign l_8[1]    = ( l_9 [1] & !i[1724]);
assign l_8[2]    = ( l_9 [2] & !i[1724]);
assign l_8[3]    = ( l_9 [3] & !i[1724]);
assign l_8[4]    = ( l_9 [4] & !i[1724]);
assign l_8[5]    = ( l_9 [5] & !i[1724]);
assign l_8[6]    = ( l_9 [6] & !i[1724]);
assign l_8[7]    = ( l_9 [7] & !i[1724]);
assign l_8[8]    = ( l_9 [8] & !i[1724]);
assign l_8[9]    = ( l_9 [9] & !i[1724]);
assign l_8[10]    = ( l_9 [10] & !i[1724]) | (      i[1724]);
assign l_8[11]    = ( l_9 [11] & !i[1724]) | (      i[1724]);
assign l_8[12]    = ( l_9 [12] & !i[1724]) | (      i[1724]);
assign l_8[13]    = ( l_9 [13] & !i[1724]) | (      i[1724]);
assign l_8[14]    = ( l_9 [14] & !i[1724]) | (      i[1724]);
assign l_8[15]    = ( l_9 [15] & !i[1724]) | (      i[1724]);
assign l_8[16]    = (!l_9 [5] & !i[1724]) | (      i[1724]);
assign l_8[17]    = ( l_9 [16] & !i[1724]) | (      i[1724]);
assign l_8[18]    = ( l_9 [17] & !i[1724]) | (      i[1724]);
assign l_8[19]    = (!l_9 [6] & !i[1724]) | (      i[1724]);
assign l_9[0]    = ( l_10 [0] & !i[1721]);
assign l_9[1]    = ( l_10 [1] & !i[1721]);
assign l_9[2]    = ( l_10 [2] & !i[1721]);
assign l_9[3]    = ( l_10 [3] & !i[1721]);
assign l_9[4]    = ( l_10 [4] & !i[1721]);
assign l_9[5]    = ( l_10 [5] & !i[1721]);
assign l_9[6]    = ( l_10 [6] & !i[1721]);
assign l_9[7]    = ( l_10 [7] & !i[1721]);
assign l_9[8]    = ( l_10 [8] & !i[1721]);
assign l_9[9]    = ( l_10 [9] & !i[1721]);
assign l_9[10]    = ( l_10 [10] & !i[1721]) | (      i[1721]);
assign l_9[11]    = ( l_10 [11] & !i[1721]) | (      i[1721]);
assign l_9[12]    = ( l_10 [12] & !i[1721]) | (      i[1721]);
assign l_9[13]    = ( l_10 [13] & !i[1721]) | (      i[1721]);
assign l_9[14]    = ( l_10 [14] & !i[1721]) | (      i[1721]);
assign l_9[15]    = ( l_10 [15] & !i[1721]) | (      i[1721]);
assign l_9[16]    = ( l_10 [16] & !i[1721]) | (      i[1721]);
assign l_9[17]    = ( l_10 [17] & !i[1721]) | (      i[1721]);

endmodule
