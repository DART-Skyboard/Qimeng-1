//circuit accuracy = 1
//test amounts  = 1000000
//total BDD nodes = 97
//total split modes = 85
//train time = 92.2647
module module_output_bit_84(i,o);

input [1893:0] i;
output  o;

wire [0:0] l_0;
wire [1:0] l_1;
wire [3:0] l_2;
wire [4:0] l_3;
wire [4:0] l_4;
wire [4:0] l_5;
wire [4:0] l_6;
wire [4:0] l_7;
wire [4:0] l_8;
wire [4:0] l_9;
wire [4:0] l_10;
wire [4:0] l_11;
wire [4:0] l_12;
wire [3:0] l_13;
wire [6:0] l_14;
wire [6:0] l_15;
wire [4:0] l_16;
wire [5:0] l_17;
wire [3:0] l_18;
wire [2:0] l_19;
wire [1:0] l_20;
wire [0:0] l_21;
wire [0:0] l_22;
wire [-1:0] l_23;

assign o = l_0[0];

assign l_0[0]    = ( l_1 [0] & !i[84]) | ( l_1 [1] &  i[84]);
assign l_1[0]    = ( l_2 [0] & !i[1722]) | ( l_2 [1] &  i[1722]);
assign l_1[1]    = ( l_2 [2] & !i[1722]) | ( l_2 [3] &  i[1722]);
assign l_2[0]    = ( l_3 [0] & !i[1723]);
assign l_2[1]    = ( l_3 [1] & !i[1723]);
assign l_2[2]    = ( l_3 [2] & !i[1723]) | (      i[1723]);
assign l_2[3]    = ( l_3 [3] & !i[1723]) | ( l_3 [4] &  i[1723]);
assign l_3[0]    = ( l_4 [0] & !i[1725]);
assign l_3[1]    = ( l_4 [1] &  i[1725]);
assign l_3[2]    = ( l_4 [2] & !i[1725]) | (      i[1725]);
assign l_3[3]    = (!i[1725]) | ( l_4 [3] &  i[1725]);
assign l_3[4]    = (!i[1725]) | ( l_4 [4] &  i[1725]);
assign l_4[0]    = ( l_5 [0] & !i[1721]);
assign l_4[1]    = ( l_5 [1] & !i[1721]);
assign l_4[2]    = ( l_5 [2] & !i[1721]) | (      i[1721]);
assign l_4[3]    = ( l_5 [3] & !i[1721]) | (      i[1721]);
assign l_4[4]    = ( l_5 [4] & !i[1721]) | (      i[1721]);
assign l_5[0]    = ( l_6 [0] & !i[1716]);
assign l_5[1]    = ( l_6 [1] & !i[1716]);
assign l_5[2]    = ( l_6 [2] & !i[1716]) | (      i[1716]);
assign l_5[3]    = ( l_6 [3] & !i[1716]) | (      i[1716]);
assign l_5[4]    = ( l_6 [4] & !i[1716]) | (      i[1716]);
assign l_6[0]    = ( l_7 [0] & !i[1717]);
assign l_6[1]    = ( l_7 [1] & !i[1717]);
assign l_6[2]    = ( l_7 [2] & !i[1717]) | (      i[1717]);
assign l_6[3]    = ( l_7 [3] & !i[1717]) | (      i[1717]);
assign l_6[4]    = ( l_7 [4] & !i[1717]) | (      i[1717]);
assign l_7[0]    = ( l_8 [0] & !i[1718]);
assign l_7[1]    = ( l_8 [1] & !i[1718]);
assign l_7[2]    = ( l_8 [2] & !i[1718]) | (      i[1718]);
assign l_7[3]    = ( l_8 [3] & !i[1718]) | (      i[1718]);
assign l_7[4]    = ( l_8 [4] & !i[1718]) | (      i[1718]);
assign l_8[0]    = ( l_9 [0] &  i[1719]);
assign l_8[1]    = ( l_9 [1] &  i[1719]);
assign l_8[2]    = (!i[1719]) | ( l_9 [2] &  i[1719]);
assign l_8[3]    = (!i[1719]) | ( l_9 [3] &  i[1719]);
assign l_8[4]    = (!i[1719]) | ( l_9 [4] &  i[1719]);
assign l_9[0]    = ( l_10 [0] & !i[1720]);
assign l_9[1]    = ( l_10 [1] & !i[1720]);
assign l_9[2]    = ( l_10 [2] & !i[1720]) | (      i[1720]);
assign l_9[3]    = ( l_10 [3] & !i[1720]) | (      i[1720]);
assign l_9[4]    = ( l_10 [4] & !i[1720]) | (      i[1720]);
assign l_10[0]    = ( l_11 [0] & !i[1724]);
assign l_10[1]    = ( l_11 [1] &  i[1724]);
assign l_10[2]    = ( l_11 [2] & !i[1724]) | (      i[1724]);
assign l_10[3]    = (!i[1724]) | ( l_11 [3] &  i[1724]);
assign l_10[4]    = ( l_11 [4] & !i[1724]) | (      i[1724]);
assign l_11[0]    = ( l_12 [0] &  i[1726]);
assign l_11[1]    = ( l_12 [1] &  i[1726]);
assign l_11[2]    = (!i[1726]) | ( l_12 [2] &  i[1726]);
assign l_11[3]    = (!i[1726]) | ( l_12 [3] &  i[1726]);
assign l_11[4]    = (!i[1726]) | ( l_12 [4] &  i[1726]);
assign l_12[0]    = ( l_13 [0] &  i[1727]);
assign l_12[1]    = ( l_13 [1] &  i[1727]);
assign l_12[2]    = (!i[1727]) | ( l_13 [2] &  i[1727]);
assign l_12[3]    = (!i[1727]) | ( l_13 [3] &  i[1727]);
assign l_12[4]    = !i[1727];
assign l_13[0]    = ( l_14 [0] & !i[1780]) | ( l_14 [1] &  i[1780]);
assign l_13[1]    = ( l_14 [2] &  i[1780]);
assign l_13[2]    = ( l_14 [3] & !i[1780]) | ( l_14 [4] &  i[1780]);
assign l_13[3]    = ( l_14 [5] & !i[1780]) | ( l_14 [6] &  i[1780]);
assign l_14[0]    = ( l_15 [0] & !i[1714]);
assign l_14[1]    = ( l_15 [1] & !i[1714]) | ( l_15 [2] &  i[1714]);
assign l_14[2]    = ( l_15 [3]);
assign l_14[3]    = ( l_15 [0] & !i[1714]) | ( l_15 [4] &  i[1714]);
assign l_14[4]    = ( l_15 [1] & !i[1714]) | (      i[1714]);
assign l_14[5]    = ( l_15 [5]);
assign l_14[6]    = ( l_15 [6]);
assign l_15[0]    = ( l_16 [0] & !i[1715]);
assign l_15[1]    = ( l_16 [0] & !i[1715]) | (      i[1715]);
assign l_15[2]    = ( l_16 [1] & !i[1715]);
assign l_15[3]    = ( l_16 [2]);
assign l_15[4]    = (!l_16 [1] & !i[1715]) | (      i[1715]);
assign l_15[5]    = ( l_16 [3]);
assign l_15[6]    = ( l_16 [4]);
assign l_16[0]    = ( l_17 [0]);
assign l_16[1]    = ( l_17 [1]);
assign l_16[2]    = ( l_17 [2] & !i[1699]) | ( l_17 [3] &  i[1699]);
assign l_16[3]    = (!l_17 [2] & !i[1699]) | ( l_17 [4] &  i[1699]);
assign l_16[4]    = (!i[1699]) | ( l_17 [5] &  i[1699]);
assign l_17[0]    = ( l_18 [0]);
assign l_17[1]    = ( l_18 [1]);
assign l_17[2]    = (!i[1700]) | ( l_18 [2] &  i[1700]);
assign l_17[3]    = ( l_18 [2] & !i[1700]);
assign l_17[4]    = (!l_18 [2] & !i[1700]) | ( l_18 [3] &  i[1700]);
assign l_17[5]    = (!i[1700]) | ( l_18 [3] &  i[1700]);
assign l_18[0]    = ( l_19 [0] & !i[1713]);
assign l_18[1]    = !i[1713];
assign l_18[2]    = ( l_19 [1]);
assign l_18[3]    = (!l_19 [1] & !i[1713]) | ( l_19 [2] &  i[1713]);
assign l_19[0]    =  i[1784];
assign l_19[1]    = ( l_20 [0]);
assign l_19[2]    = (!l_20 [0] & !i[1784]) | ( l_20 [1] &  i[1784]);
assign l_20[0]    = ( l_21 [0] & !i[1696]);
assign l_20[1]    = (!l_21 [0] & !i[1696]) | (      i[1696]);
assign l_21[0]    = ( l_22 [0] & !i[1697]);
assign l_22[0]    = !i[1698];

endmodule
