module RISCV_train(input_data_all, output_data_all);

input	[1796:0]	input_data_all;
wire	[1825:0]	output_data_all;

module_output_bit_0	m0	(input_data_all[1796:0],output_data_all[0]);
module_output_bit_1	m1	(input_data_all[1796:0],output_data_all[1]);
module_output_bit_2	m2	(input_data_all[1796:0],output_data_all[2]);
module_output_bit_3	m3	(input_data_all[1796:0],output_data_all[3]);
module_output_bit_4	m4	(input_data_all[1796:0],output_data_all[4]);
module_output_bit_5	m5	(input_data_all[1796:0],output_data_all[5]);
module_output_bit_6	m6	(input_data_all[1796:0],output_data_all[6]);
module_output_bit_7	m7	(input_data_all[1796:0],output_data_all[7]);
module_output_bit_8	m8	(input_data_all[1796:0],output_data_all[8]);
module_output_bit_9	m9	(input_data_all[1796:0],output_data_all[9]);
module_output_bit_10	m10	(input_data_all[1796:0],output_data_all[10]);
module_output_bit_11	m11	(input_data_all[1796:0],output_data_all[11]);
module_output_bit_12	m12	(input_data_all[1796:0],output_data_all[12]);
module_output_bit_13	m13	(input_data_all[1796:0],output_data_all[13]);
module_output_bit_14	m14	(input_data_all[1796:0],output_data_all[14]);
module_output_bit_15	m15	(input_data_all[1796:0],output_data_all[15]);
module_output_bit_16	m16	(input_data_all[1796:0],output_data_all[16]);
module_output_bit_17	m17	(input_data_all[1796:0],output_data_all[17]);
module_output_bit_18	m18	(input_data_all[1796:0],output_data_all[18]);
module_output_bit_19	m19	(input_data_all[1796:0],output_data_all[19]);
module_output_bit_20	m20	(input_data_all[1796:0],output_data_all[20]);
module_output_bit_21	m21	(input_data_all[1796:0],output_data_all[21]);
module_output_bit_22	m22	(input_data_all[1796:0],output_data_all[22]);
module_output_bit_23	m23	(input_data_all[1796:0],output_data_all[23]);
module_output_bit_24	m24	(input_data_all[1796:0],output_data_all[24]);
module_output_bit_25	m25	(input_data_all[1796:0],output_data_all[25]);
module_output_bit_26	m26	(input_data_all[1796:0],output_data_all[26]);
module_output_bit_27	m27	(input_data_all[1796:0],output_data_all[27]);
module_output_bit_28	m28	(input_data_all[1796:0],output_data_all[28]);
module_output_bit_29	m29	(input_data_all[1796:0],output_data_all[29]);
module_output_bit_30	m30	(input_data_all[1796:0],output_data_all[30]);
module_output_bit_31	m31	(input_data_all[1796:0],output_data_all[31]);
module_output_bit_32	m32	(input_data_all[1796:0],output_data_all[32]);
module_output_bit_33	m33	(input_data_all[1796:0],output_data_all[33]);
module_output_bit_34	m34	(input_data_all[1796:0],output_data_all[34]);
module_output_bit_35	m35	(input_data_all[1796:0],output_data_all[35]);
module_output_bit_36	m36	(input_data_all[1796:0],output_data_all[36]);
module_output_bit_37	m37	(input_data_all[1796:0],output_data_all[37]);
module_output_bit_38	m38	(input_data_all[1796:0],output_data_all[38]);
module_output_bit_39	m39	(input_data_all[1796:0],output_data_all[39]);
module_output_bit_40	m40	(input_data_all[1796:0],output_data_all[40]);
module_output_bit_41	m41	(input_data_all[1796:0],output_data_all[41]);
module_output_bit_42	m42	(input_data_all[1796:0],output_data_all[42]);
module_output_bit_43	m43	(input_data_all[1796:0],output_data_all[43]);
module_output_bit_44	m44	(input_data_all[1796:0],output_data_all[44]);
module_output_bit_45	m45	(input_data_all[1796:0],output_data_all[45]);
module_output_bit_46	m46	(input_data_all[1796:0],output_data_all[46]);
module_output_bit_47	m47	(input_data_all[1796:0],output_data_all[47]);
module_output_bit_48	m48	(input_data_all[1796:0],output_data_all[48]);
module_output_bit_49	m49	(input_data_all[1796:0],output_data_all[49]);
module_output_bit_50	m50	(input_data_all[1796:0],output_data_all[50]);
module_output_bit_51	m51	(input_data_all[1796:0],output_data_all[51]);
module_output_bit_52	m52	(input_data_all[1796:0],output_data_all[52]);
module_output_bit_53	m53	(input_data_all[1796:0],output_data_all[53]);
module_output_bit_54	m54	(input_data_all[1796:0],output_data_all[54]);
module_output_bit_55	m55	(input_data_all[1796:0],output_data_all[55]);
module_output_bit_56	m56	(input_data_all[1796:0],output_data_all[56]);
module_output_bit_57	m57	(input_data_all[1796:0],output_data_all[57]);
module_output_bit_58	m58	(input_data_all[1796:0],output_data_all[58]);
module_output_bit_59	m59	(input_data_all[1796:0],output_data_all[59]);
module_output_bit_60	m60	(input_data_all[1796:0],output_data_all[60]);
module_output_bit_61	m61	(input_data_all[1796:0],output_data_all[61]);
module_output_bit_62	m62	(input_data_all[1796:0],output_data_all[62]);
module_output_bit_63	m63	(input_data_all[1796:0],output_data_all[63]);
module_output_bit_64	m64	(input_data_all[1796:0],output_data_all[64]);
module_output_bit_65	m65	(input_data_all[1796:0],output_data_all[65]);
module_output_bit_66	m66	(input_data_all[1796:0],output_data_all[66]);
module_output_bit_67	m67	(input_data_all[1796:0],output_data_all[67]);
module_output_bit_68	m68	(input_data_all[1796:0],output_data_all[68]);
module_output_bit_69	m69	(input_data_all[1796:0],output_data_all[69]);
module_output_bit_70	m70	(input_data_all[1796:0],output_data_all[70]);
module_output_bit_71	m71	(input_data_all[1796:0],output_data_all[71]);
module_output_bit_72	m72	(input_data_all[1796:0],output_data_all[72]);
module_output_bit_73	m73	(input_data_all[1796:0],output_data_all[73]);
module_output_bit_74	m74	(input_data_all[1796:0],output_data_all[74]);
module_output_bit_75	m75	(input_data_all[1796:0],output_data_all[75]);
module_output_bit_76	m76	(input_data_all[1796:0],output_data_all[76]);
module_output_bit_77	m77	(input_data_all[1796:0],output_data_all[77]);
module_output_bit_78	m78	(input_data_all[1796:0],output_data_all[78]);
module_output_bit_79	m79	(input_data_all[1796:0],output_data_all[79]);
module_output_bit_80	m80	(input_data_all[1796:0],output_data_all[80]);
module_output_bit_81	m81	(input_data_all[1796:0],output_data_all[81]);
module_output_bit_82	m82	(input_data_all[1796:0],output_data_all[82]);
module_output_bit_83	m83	(input_data_all[1796:0],output_data_all[83]);
module_output_bit_84	m84	(input_data_all[1796:0],output_data_all[84]);
module_output_bit_85	m85	(input_data_all[1796:0],output_data_all[85]);
module_output_bit_86	m86	(input_data_all[1796:0],output_data_all[86]);
module_output_bit_87	m87	(input_data_all[1796:0],output_data_all[87]);
module_output_bit_88	m88	(input_data_all[1796:0],output_data_all[88]);
module_output_bit_89	m89	(input_data_all[1796:0],output_data_all[89]);
module_output_bit_90	m90	(input_data_all[1796:0],output_data_all[90]);
module_output_bit_91	m91	(input_data_all[1796:0],output_data_all[91]);
module_output_bit_92	m92	(input_data_all[1796:0],output_data_all[92]);
module_output_bit_93	m93	(input_data_all[1796:0],output_data_all[93]);
module_output_bit_94	m94	(input_data_all[1796:0],output_data_all[94]);
module_output_bit_95	m95	(input_data_all[1796:0],output_data_all[95]);
module_output_bit_96	m96	(input_data_all[1796:0],output_data_all[96]);
module_output_bit_97	m97	(input_data_all[1796:0],output_data_all[97]);
module_output_bit_98	m98	(input_data_all[1796:0],output_data_all[98]);
module_output_bit_99	m99	(input_data_all[1796:0],output_data_all[99]);
module_output_bit_100	m100	(input_data_all[1796:0],output_data_all[100]);
module_output_bit_101	m101	(input_data_all[1796:0],output_data_all[101]);
module_output_bit_102	m102	(input_data_all[1796:0],output_data_all[102]);
module_output_bit_103	m103	(input_data_all[1796:0],output_data_all[103]);
module_output_bit_104	m104	(input_data_all[1796:0],output_data_all[104]);
module_output_bit_105	m105	(input_data_all[1796:0],output_data_all[105]);
module_output_bit_106	m106	(input_data_all[1796:0],output_data_all[106]);
module_output_bit_107	m107	(input_data_all[1796:0],output_data_all[107]);
module_output_bit_108	m108	(input_data_all[1796:0],output_data_all[108]);
module_output_bit_109	m109	(input_data_all[1796:0],output_data_all[109]);
module_output_bit_110	m110	(input_data_all[1796:0],output_data_all[110]);
module_output_bit_111	m111	(input_data_all[1796:0],output_data_all[111]);
module_output_bit_112	m112	(input_data_all[1796:0],output_data_all[112]);
module_output_bit_113	m113	(input_data_all[1796:0],output_data_all[113]);
module_output_bit_114	m114	(input_data_all[1796:0],output_data_all[114]);
module_output_bit_115	m115	(input_data_all[1796:0],output_data_all[115]);
module_output_bit_116	m116	(input_data_all[1796:0],output_data_all[116]);
module_output_bit_117	m117	(input_data_all[1796:0],output_data_all[117]);
module_output_bit_118	m118	(input_data_all[1796:0],output_data_all[118]);
module_output_bit_119	m119	(input_data_all[1796:0],output_data_all[119]);
module_output_bit_120	m120	(input_data_all[1796:0],output_data_all[120]);
module_output_bit_121	m121	(input_data_all[1796:0],output_data_all[121]);
module_output_bit_122	m122	(input_data_all[1796:0],output_data_all[122]);
module_output_bit_123	m123	(input_data_all[1796:0],output_data_all[123]);
module_output_bit_124	m124	(input_data_all[1796:0],output_data_all[124]);
module_output_bit_125	m125	(input_data_all[1796:0],output_data_all[125]);
module_output_bit_126	m126	(input_data_all[1796:0],output_data_all[126]);
module_output_bit_127	m127	(input_data_all[1796:0],output_data_all[127]);
module_output_bit_128	m128	(input_data_all[1796:0],output_data_all[128]);
module_output_bit_129	m129	(input_data_all[1796:0],output_data_all[129]);
module_output_bit_130	m130	(input_data_all[1796:0],output_data_all[130]);
module_output_bit_131	m131	(input_data_all[1796:0],output_data_all[131]);
module_output_bit_132	m132	(input_data_all[1796:0],output_data_all[132]);
module_output_bit_133	m133	(input_data_all[1796:0],output_data_all[133]);
module_output_bit_134	m134	(input_data_all[1796:0],output_data_all[134]);
module_output_bit_135	m135	(input_data_all[1796:0],output_data_all[135]);
module_output_bit_136	m136	(input_data_all[1796:0],output_data_all[136]);
module_output_bit_137	m137	(input_data_all[1796:0],output_data_all[137]);
module_output_bit_138	m138	(input_data_all[1796:0],output_data_all[138]);
module_output_bit_139	m139	(input_data_all[1796:0],output_data_all[139]);
module_output_bit_140	m140	(input_data_all[1796:0],output_data_all[140]);
module_output_bit_141	m141	(input_data_all[1796:0],output_data_all[141]);
module_output_bit_142	m142	(input_data_all[1796:0],output_data_all[142]);
module_output_bit_143	m143	(input_data_all[1796:0],output_data_all[143]);
module_output_bit_144	m144	(input_data_all[1796:0],output_data_all[144]);
module_output_bit_145	m145	(input_data_all[1796:0],output_data_all[145]);
module_output_bit_146	m146	(input_data_all[1796:0],output_data_all[146]);
module_output_bit_147	m147	(input_data_all[1796:0],output_data_all[147]);
module_output_bit_148	m148	(input_data_all[1796:0],output_data_all[148]);
module_output_bit_149	m149	(input_data_all[1796:0],output_data_all[149]);
module_output_bit_150	m150	(input_data_all[1796:0],output_data_all[150]);
module_output_bit_151	m151	(input_data_all[1796:0],output_data_all[151]);
module_output_bit_152	m152	(input_data_all[1796:0],output_data_all[152]);
module_output_bit_153	m153	(input_data_all[1796:0],output_data_all[153]);
module_output_bit_154	m154	(input_data_all[1796:0],output_data_all[154]);
module_output_bit_155	m155	(input_data_all[1796:0],output_data_all[155]);
module_output_bit_156	m156	(input_data_all[1796:0],output_data_all[156]);
module_output_bit_157	m157	(input_data_all[1796:0],output_data_all[157]);
module_output_bit_158	m158	(input_data_all[1796:0],output_data_all[158]);
module_output_bit_159	m159	(input_data_all[1796:0],output_data_all[159]);
module_output_bit_160	m160	(input_data_all[1796:0],output_data_all[160]);
module_output_bit_161	m161	(input_data_all[1796:0],output_data_all[161]);
module_output_bit_162	m162	(input_data_all[1796:0],output_data_all[162]);
module_output_bit_163	m163	(input_data_all[1796:0],output_data_all[163]);
module_output_bit_164	m164	(input_data_all[1796:0],output_data_all[164]);
module_output_bit_165	m165	(input_data_all[1796:0],output_data_all[165]);
module_output_bit_166	m166	(input_data_all[1796:0],output_data_all[166]);
module_output_bit_167	m167	(input_data_all[1796:0],output_data_all[167]);
module_output_bit_168	m168	(input_data_all[1796:0],output_data_all[168]);
module_output_bit_169	m169	(input_data_all[1796:0],output_data_all[169]);
module_output_bit_170	m170	(input_data_all[1796:0],output_data_all[170]);
module_output_bit_171	m171	(input_data_all[1796:0],output_data_all[171]);
module_output_bit_172	m172	(input_data_all[1796:0],output_data_all[172]);
module_output_bit_173	m173	(input_data_all[1796:0],output_data_all[173]);
module_output_bit_174	m174	(input_data_all[1796:0],output_data_all[174]);
module_output_bit_175	m175	(input_data_all[1796:0],output_data_all[175]);
module_output_bit_176	m176	(input_data_all[1796:0],output_data_all[176]);
module_output_bit_177	m177	(input_data_all[1796:0],output_data_all[177]);
module_output_bit_178	m178	(input_data_all[1796:0],output_data_all[178]);
module_output_bit_179	m179	(input_data_all[1796:0],output_data_all[179]);
module_output_bit_180	m180	(input_data_all[1796:0],output_data_all[180]);
module_output_bit_181	m181	(input_data_all[1796:0],output_data_all[181]);
module_output_bit_182	m182	(input_data_all[1796:0],output_data_all[182]);
module_output_bit_183	m183	(input_data_all[1796:0],output_data_all[183]);
module_output_bit_184	m184	(input_data_all[1796:0],output_data_all[184]);
module_output_bit_185	m185	(input_data_all[1796:0],output_data_all[185]);
module_output_bit_186	m186	(input_data_all[1796:0],output_data_all[186]);
module_output_bit_187	m187	(input_data_all[1796:0],output_data_all[187]);
module_output_bit_188	m188	(input_data_all[1796:0],output_data_all[188]);
module_output_bit_189	m189	(input_data_all[1796:0],output_data_all[189]);
module_output_bit_190	m190	(input_data_all[1796:0],output_data_all[190]);
module_output_bit_191	m191	(input_data_all[1796:0],output_data_all[191]);
module_output_bit_192	m192	(input_data_all[1796:0],output_data_all[192]);
module_output_bit_193	m193	(input_data_all[1796:0],output_data_all[193]);
module_output_bit_194	m194	(input_data_all[1796:0],output_data_all[194]);
module_output_bit_195	m195	(input_data_all[1796:0],output_data_all[195]);
module_output_bit_196	m196	(input_data_all[1796:0],output_data_all[196]);
module_output_bit_197	m197	(input_data_all[1796:0],output_data_all[197]);
module_output_bit_198	m198	(input_data_all[1796:0],output_data_all[198]);
module_output_bit_199	m199	(input_data_all[1796:0],output_data_all[199]);
module_output_bit_200	m200	(input_data_all[1796:0],output_data_all[200]);
module_output_bit_201	m201	(input_data_all[1796:0],output_data_all[201]);
module_output_bit_202	m202	(input_data_all[1796:0],output_data_all[202]);
module_output_bit_203	m203	(input_data_all[1796:0],output_data_all[203]);
module_output_bit_204	m204	(input_data_all[1796:0],output_data_all[204]);
module_output_bit_205	m205	(input_data_all[1796:0],output_data_all[205]);
module_output_bit_206	m206	(input_data_all[1796:0],output_data_all[206]);
module_output_bit_207	m207	(input_data_all[1796:0],output_data_all[207]);
module_output_bit_208	m208	(input_data_all[1796:0],output_data_all[208]);
module_output_bit_209	m209	(input_data_all[1796:0],output_data_all[209]);
module_output_bit_210	m210	(input_data_all[1796:0],output_data_all[210]);
module_output_bit_211	m211	(input_data_all[1796:0],output_data_all[211]);
module_output_bit_212	m212	(input_data_all[1796:0],output_data_all[212]);
module_output_bit_213	m213	(input_data_all[1796:0],output_data_all[213]);
module_output_bit_214	m214	(input_data_all[1796:0],output_data_all[214]);
module_output_bit_215	m215	(input_data_all[1796:0],output_data_all[215]);
module_output_bit_216	m216	(input_data_all[1796:0],output_data_all[216]);
module_output_bit_217	m217	(input_data_all[1796:0],output_data_all[217]);
module_output_bit_218	m218	(input_data_all[1796:0],output_data_all[218]);
module_output_bit_219	m219	(input_data_all[1796:0],output_data_all[219]);
module_output_bit_220	m220	(input_data_all[1796:0],output_data_all[220]);
module_output_bit_221	m221	(input_data_all[1796:0],output_data_all[221]);
module_output_bit_222	m222	(input_data_all[1796:0],output_data_all[222]);
module_output_bit_223	m223	(input_data_all[1796:0],output_data_all[223]);
module_output_bit_224	m224	(input_data_all[1796:0],output_data_all[224]);
module_output_bit_225	m225	(input_data_all[1796:0],output_data_all[225]);
module_output_bit_226	m226	(input_data_all[1796:0],output_data_all[226]);
module_output_bit_227	m227	(input_data_all[1796:0],output_data_all[227]);
module_output_bit_228	m228	(input_data_all[1796:0],output_data_all[228]);
module_output_bit_229	m229	(input_data_all[1796:0],output_data_all[229]);
module_output_bit_230	m230	(input_data_all[1796:0],output_data_all[230]);
module_output_bit_231	m231	(input_data_all[1796:0],output_data_all[231]);
module_output_bit_232	m232	(input_data_all[1796:0],output_data_all[232]);
module_output_bit_233	m233	(input_data_all[1796:0],output_data_all[233]);
module_output_bit_234	m234	(input_data_all[1796:0],output_data_all[234]);
module_output_bit_235	m235	(input_data_all[1796:0],output_data_all[235]);
module_output_bit_236	m236	(input_data_all[1796:0],output_data_all[236]);
module_output_bit_237	m237	(input_data_all[1796:0],output_data_all[237]);
module_output_bit_238	m238	(input_data_all[1796:0],output_data_all[238]);
module_output_bit_239	m239	(input_data_all[1796:0],output_data_all[239]);
module_output_bit_240	m240	(input_data_all[1796:0],output_data_all[240]);
module_output_bit_241	m241	(input_data_all[1796:0],output_data_all[241]);
module_output_bit_242	m242	(input_data_all[1796:0],output_data_all[242]);
module_output_bit_243	m243	(input_data_all[1796:0],output_data_all[243]);
module_output_bit_244	m244	(input_data_all[1796:0],output_data_all[244]);
module_output_bit_245	m245	(input_data_all[1796:0],output_data_all[245]);
module_output_bit_246	m246	(input_data_all[1796:0],output_data_all[246]);
module_output_bit_247	m247	(input_data_all[1796:0],output_data_all[247]);
module_output_bit_248	m248	(input_data_all[1796:0],output_data_all[248]);
module_output_bit_249	m249	(input_data_all[1796:0],output_data_all[249]);
module_output_bit_250	m250	(input_data_all[1796:0],output_data_all[250]);
module_output_bit_251	m251	(input_data_all[1796:0],output_data_all[251]);
module_output_bit_252	m252	(input_data_all[1796:0],output_data_all[252]);
module_output_bit_253	m253	(input_data_all[1796:0],output_data_all[253]);
module_output_bit_254	m254	(input_data_all[1796:0],output_data_all[254]);
module_output_bit_255	m255	(input_data_all[1796:0],output_data_all[255]);
module_output_bit_256	m256	(input_data_all[1796:0],output_data_all[256]);
module_output_bit_257	m257	(input_data_all[1796:0],output_data_all[257]);
module_output_bit_258	m258	(input_data_all[1796:0],output_data_all[258]);
module_output_bit_259	m259	(input_data_all[1796:0],output_data_all[259]);
module_output_bit_260	m260	(input_data_all[1796:0],output_data_all[260]);
module_output_bit_261	m261	(input_data_all[1796:0],output_data_all[261]);
module_output_bit_262	m262	(input_data_all[1796:0],output_data_all[262]);
module_output_bit_263	m263	(input_data_all[1796:0],output_data_all[263]);
module_output_bit_264	m264	(input_data_all[1796:0],output_data_all[264]);
module_output_bit_265	m265	(input_data_all[1796:0],output_data_all[265]);
module_output_bit_266	m266	(input_data_all[1796:0],output_data_all[266]);
module_output_bit_267	m267	(input_data_all[1796:0],output_data_all[267]);
module_output_bit_268	m268	(input_data_all[1796:0],output_data_all[268]);
module_output_bit_269	m269	(input_data_all[1796:0],output_data_all[269]);
module_output_bit_270	m270	(input_data_all[1796:0],output_data_all[270]);
module_output_bit_271	m271	(input_data_all[1796:0],output_data_all[271]);
module_output_bit_272	m272	(input_data_all[1796:0],output_data_all[272]);
module_output_bit_273	m273	(input_data_all[1796:0],output_data_all[273]);
module_output_bit_274	m274	(input_data_all[1796:0],output_data_all[274]);
module_output_bit_275	m275	(input_data_all[1796:0],output_data_all[275]);
module_output_bit_276	m276	(input_data_all[1796:0],output_data_all[276]);
module_output_bit_277	m277	(input_data_all[1796:0],output_data_all[277]);
module_output_bit_278	m278	(input_data_all[1796:0],output_data_all[278]);
module_output_bit_279	m279	(input_data_all[1796:0],output_data_all[279]);
module_output_bit_280	m280	(input_data_all[1796:0],output_data_all[280]);
module_output_bit_281	m281	(input_data_all[1796:0],output_data_all[281]);
module_output_bit_282	m282	(input_data_all[1796:0],output_data_all[282]);
module_output_bit_283	m283	(input_data_all[1796:0],output_data_all[283]);
module_output_bit_284	m284	(input_data_all[1796:0],output_data_all[284]);
module_output_bit_285	m285	(input_data_all[1796:0],output_data_all[285]);
module_output_bit_286	m286	(input_data_all[1796:0],output_data_all[286]);
module_output_bit_287	m287	(input_data_all[1796:0],output_data_all[287]);
module_output_bit_288	m288	(input_data_all[1796:0],output_data_all[288]);
module_output_bit_289	m289	(input_data_all[1796:0],output_data_all[289]);
module_output_bit_290	m290	(input_data_all[1796:0],output_data_all[290]);
module_output_bit_291	m291	(input_data_all[1796:0],output_data_all[291]);
module_output_bit_292	m292	(input_data_all[1796:0],output_data_all[292]);
module_output_bit_293	m293	(input_data_all[1796:0],output_data_all[293]);
module_output_bit_294	m294	(input_data_all[1796:0],output_data_all[294]);
module_output_bit_295	m295	(input_data_all[1796:0],output_data_all[295]);
module_output_bit_296	m296	(input_data_all[1796:0],output_data_all[296]);
module_output_bit_297	m297	(input_data_all[1796:0],output_data_all[297]);
module_output_bit_298	m298	(input_data_all[1796:0],output_data_all[298]);
module_output_bit_299	m299	(input_data_all[1796:0],output_data_all[299]);
module_output_bit_300	m300	(input_data_all[1796:0],output_data_all[300]);
module_output_bit_301	m301	(input_data_all[1796:0],output_data_all[301]);
module_output_bit_302	m302	(input_data_all[1796:0],output_data_all[302]);
module_output_bit_303	m303	(input_data_all[1796:0],output_data_all[303]);
module_output_bit_304	m304	(input_data_all[1796:0],output_data_all[304]);
module_output_bit_305	m305	(input_data_all[1796:0],output_data_all[305]);
module_output_bit_306	m306	(input_data_all[1796:0],output_data_all[306]);
module_output_bit_307	m307	(input_data_all[1796:0],output_data_all[307]);
module_output_bit_308	m308	(input_data_all[1796:0],output_data_all[308]);
module_output_bit_309	m309	(input_data_all[1796:0],output_data_all[309]);
module_output_bit_310	m310	(input_data_all[1796:0],output_data_all[310]);
module_output_bit_311	m311	(input_data_all[1796:0],output_data_all[311]);
module_output_bit_312	m312	(input_data_all[1796:0],output_data_all[312]);
module_output_bit_313	m313	(input_data_all[1796:0],output_data_all[313]);
module_output_bit_314	m314	(input_data_all[1796:0],output_data_all[314]);
module_output_bit_315	m315	(input_data_all[1796:0],output_data_all[315]);
module_output_bit_316	m316	(input_data_all[1796:0],output_data_all[316]);
module_output_bit_317	m317	(input_data_all[1796:0],output_data_all[317]);
module_output_bit_318	m318	(input_data_all[1796:0],output_data_all[318]);
module_output_bit_319	m319	(input_data_all[1796:0],output_data_all[319]);
module_output_bit_320	m320	(input_data_all[1796:0],output_data_all[320]);
module_output_bit_321	m321	(input_data_all[1796:0],output_data_all[321]);
module_output_bit_322	m322	(input_data_all[1796:0],output_data_all[322]);
module_output_bit_323	m323	(input_data_all[1796:0],output_data_all[323]);
module_output_bit_324	m324	(input_data_all[1796:0],output_data_all[324]);
module_output_bit_325	m325	(input_data_all[1796:0],output_data_all[325]);
module_output_bit_326	m326	(input_data_all[1796:0],output_data_all[326]);
module_output_bit_327	m327	(input_data_all[1796:0],output_data_all[327]);
module_output_bit_328	m328	(input_data_all[1796:0],output_data_all[328]);
module_output_bit_329	m329	(input_data_all[1796:0],output_data_all[329]);
module_output_bit_330	m330	(input_data_all[1796:0],output_data_all[330]);
module_output_bit_331	m331	(input_data_all[1796:0],output_data_all[331]);
module_output_bit_332	m332	(input_data_all[1796:0],output_data_all[332]);
module_output_bit_333	m333	(input_data_all[1796:0],output_data_all[333]);
module_output_bit_334	m334	(input_data_all[1796:0],output_data_all[334]);
module_output_bit_335	m335	(input_data_all[1796:0],output_data_all[335]);
module_output_bit_336	m336	(input_data_all[1796:0],output_data_all[336]);
module_output_bit_337	m337	(input_data_all[1796:0],output_data_all[337]);
module_output_bit_338	m338	(input_data_all[1796:0],output_data_all[338]);
module_output_bit_339	m339	(input_data_all[1796:0],output_data_all[339]);
module_output_bit_340	m340	(input_data_all[1796:0],output_data_all[340]);
module_output_bit_341	m341	(input_data_all[1796:0],output_data_all[341]);
module_output_bit_342	m342	(input_data_all[1796:0],output_data_all[342]);
module_output_bit_343	m343	(input_data_all[1796:0],output_data_all[343]);
module_output_bit_344	m344	(input_data_all[1796:0],output_data_all[344]);
module_output_bit_345	m345	(input_data_all[1796:0],output_data_all[345]);
module_output_bit_346	m346	(input_data_all[1796:0],output_data_all[346]);
module_output_bit_347	m347	(input_data_all[1796:0],output_data_all[347]);
module_output_bit_348	m348	(input_data_all[1796:0],output_data_all[348]);
module_output_bit_349	m349	(input_data_all[1796:0],output_data_all[349]);
module_output_bit_350	m350	(input_data_all[1796:0],output_data_all[350]);
module_output_bit_351	m351	(input_data_all[1796:0],output_data_all[351]);
module_output_bit_352	m352	(input_data_all[1796:0],output_data_all[352]);
module_output_bit_353	m353	(input_data_all[1796:0],output_data_all[353]);
module_output_bit_354	m354	(input_data_all[1796:0],output_data_all[354]);
module_output_bit_355	m355	(input_data_all[1796:0],output_data_all[355]);
module_output_bit_356	m356	(input_data_all[1796:0],output_data_all[356]);
module_output_bit_357	m357	(input_data_all[1796:0],output_data_all[357]);
module_output_bit_358	m358	(input_data_all[1796:0],output_data_all[358]);
module_output_bit_359	m359	(input_data_all[1796:0],output_data_all[359]);
module_output_bit_360	m360	(input_data_all[1796:0],output_data_all[360]);
module_output_bit_361	m361	(input_data_all[1796:0],output_data_all[361]);
module_output_bit_362	m362	(input_data_all[1796:0],output_data_all[362]);
module_output_bit_363	m363	(input_data_all[1796:0],output_data_all[363]);
module_output_bit_364	m364	(input_data_all[1796:0],output_data_all[364]);
module_output_bit_365	m365	(input_data_all[1796:0],output_data_all[365]);
module_output_bit_366	m366	(input_data_all[1796:0],output_data_all[366]);
module_output_bit_367	m367	(input_data_all[1796:0],output_data_all[367]);
module_output_bit_368	m368	(input_data_all[1796:0],output_data_all[368]);
module_output_bit_369	m369	(input_data_all[1796:0],output_data_all[369]);
module_output_bit_370	m370	(input_data_all[1796:0],output_data_all[370]);
module_output_bit_371	m371	(input_data_all[1796:0],output_data_all[371]);
module_output_bit_372	m372	(input_data_all[1796:0],output_data_all[372]);
module_output_bit_373	m373	(input_data_all[1796:0],output_data_all[373]);
module_output_bit_374	m374	(input_data_all[1796:0],output_data_all[374]);
module_output_bit_375	m375	(input_data_all[1796:0],output_data_all[375]);
module_output_bit_376	m376	(input_data_all[1796:0],output_data_all[376]);
module_output_bit_377	m377	(input_data_all[1796:0],output_data_all[377]);
module_output_bit_378	m378	(input_data_all[1796:0],output_data_all[378]);
module_output_bit_379	m379	(input_data_all[1796:0],output_data_all[379]);
module_output_bit_380	m380	(input_data_all[1796:0],output_data_all[380]);
module_output_bit_381	m381	(input_data_all[1796:0],output_data_all[381]);
module_output_bit_382	m382	(input_data_all[1796:0],output_data_all[382]);
module_output_bit_383	m383	(input_data_all[1796:0],output_data_all[383]);
module_output_bit_384	m384	(input_data_all[1796:0],output_data_all[384]);
module_output_bit_385	m385	(input_data_all[1796:0],output_data_all[385]);
module_output_bit_386	m386	(input_data_all[1796:0],output_data_all[386]);
module_output_bit_387	m387	(input_data_all[1796:0],output_data_all[387]);
module_output_bit_388	m388	(input_data_all[1796:0],output_data_all[388]);
module_output_bit_389	m389	(input_data_all[1796:0],output_data_all[389]);
module_output_bit_390	m390	(input_data_all[1796:0],output_data_all[390]);
module_output_bit_391	m391	(input_data_all[1796:0],output_data_all[391]);
module_output_bit_392	m392	(input_data_all[1796:0],output_data_all[392]);
module_output_bit_393	m393	(input_data_all[1796:0],output_data_all[393]);
module_output_bit_394	m394	(input_data_all[1796:0],output_data_all[394]);
module_output_bit_395	m395	(input_data_all[1796:0],output_data_all[395]);
module_output_bit_396	m396	(input_data_all[1796:0],output_data_all[396]);
module_output_bit_397	m397	(input_data_all[1796:0],output_data_all[397]);
module_output_bit_398	m398	(input_data_all[1796:0],output_data_all[398]);
module_output_bit_399	m399	(input_data_all[1796:0],output_data_all[399]);
module_output_bit_400	m400	(input_data_all[1796:0],output_data_all[400]);
module_output_bit_401	m401	(input_data_all[1796:0],output_data_all[401]);
module_output_bit_402	m402	(input_data_all[1796:0],output_data_all[402]);
module_output_bit_403	m403	(input_data_all[1796:0],output_data_all[403]);
module_output_bit_404	m404	(input_data_all[1796:0],output_data_all[404]);
module_output_bit_405	m405	(input_data_all[1796:0],output_data_all[405]);
module_output_bit_406	m406	(input_data_all[1796:0],output_data_all[406]);
module_output_bit_407	m407	(input_data_all[1796:0],output_data_all[407]);
module_output_bit_408	m408	(input_data_all[1796:0],output_data_all[408]);
module_output_bit_409	m409	(input_data_all[1796:0],output_data_all[409]);
module_output_bit_410	m410	(input_data_all[1796:0],output_data_all[410]);
module_output_bit_411	m411	(input_data_all[1796:0],output_data_all[411]);
module_output_bit_412	m412	(input_data_all[1796:0],output_data_all[412]);
module_output_bit_413	m413	(input_data_all[1796:0],output_data_all[413]);
module_output_bit_414	m414	(input_data_all[1796:0],output_data_all[414]);
module_output_bit_415	m415	(input_data_all[1796:0],output_data_all[415]);
module_output_bit_416	m416	(input_data_all[1796:0],output_data_all[416]);
module_output_bit_417	m417	(input_data_all[1796:0],output_data_all[417]);
module_output_bit_418	m418	(input_data_all[1796:0],output_data_all[418]);
module_output_bit_419	m419	(input_data_all[1796:0],output_data_all[419]);
module_output_bit_420	m420	(input_data_all[1796:0],output_data_all[420]);
module_output_bit_421	m421	(input_data_all[1796:0],output_data_all[421]);
module_output_bit_422	m422	(input_data_all[1796:0],output_data_all[422]);
module_output_bit_423	m423	(input_data_all[1796:0],output_data_all[423]);
module_output_bit_424	m424	(input_data_all[1796:0],output_data_all[424]);
module_output_bit_425	m425	(input_data_all[1796:0],output_data_all[425]);
module_output_bit_426	m426	(input_data_all[1796:0],output_data_all[426]);
module_output_bit_427	m427	(input_data_all[1796:0],output_data_all[427]);
module_output_bit_428	m428	(input_data_all[1796:0],output_data_all[428]);
module_output_bit_429	m429	(input_data_all[1796:0],output_data_all[429]);
module_output_bit_430	m430	(input_data_all[1796:0],output_data_all[430]);
module_output_bit_431	m431	(input_data_all[1796:0],output_data_all[431]);
module_output_bit_432	m432	(input_data_all[1796:0],output_data_all[432]);
module_output_bit_433	m433	(input_data_all[1796:0],output_data_all[433]);
module_output_bit_434	m434	(input_data_all[1796:0],output_data_all[434]);
module_output_bit_435	m435	(input_data_all[1796:0],output_data_all[435]);
module_output_bit_436	m436	(input_data_all[1796:0],output_data_all[436]);
module_output_bit_437	m437	(input_data_all[1796:0],output_data_all[437]);
module_output_bit_438	m438	(input_data_all[1796:0],output_data_all[438]);
module_output_bit_439	m439	(input_data_all[1796:0],output_data_all[439]);
module_output_bit_440	m440	(input_data_all[1796:0],output_data_all[440]);
module_output_bit_441	m441	(input_data_all[1796:0],output_data_all[441]);
module_output_bit_442	m442	(input_data_all[1796:0],output_data_all[442]);
module_output_bit_443	m443	(input_data_all[1796:0],output_data_all[443]);
module_output_bit_444	m444	(input_data_all[1796:0],output_data_all[444]);
module_output_bit_445	m445	(input_data_all[1796:0],output_data_all[445]);
module_output_bit_446	m446	(input_data_all[1796:0],output_data_all[446]);
module_output_bit_447	m447	(input_data_all[1796:0],output_data_all[447]);
module_output_bit_448	m448	(input_data_all[1796:0],output_data_all[448]);
module_output_bit_449	m449	(input_data_all[1796:0],output_data_all[449]);
module_output_bit_450	m450	(input_data_all[1796:0],output_data_all[450]);
module_output_bit_451	m451	(input_data_all[1796:0],output_data_all[451]);
module_output_bit_452	m452	(input_data_all[1796:0],output_data_all[452]);
module_output_bit_453	m453	(input_data_all[1796:0],output_data_all[453]);
module_output_bit_454	m454	(input_data_all[1796:0],output_data_all[454]);
module_output_bit_455	m455	(input_data_all[1796:0],output_data_all[455]);
module_output_bit_456	m456	(input_data_all[1796:0],output_data_all[456]);
module_output_bit_457	m457	(input_data_all[1796:0],output_data_all[457]);
module_output_bit_458	m458	(input_data_all[1796:0],output_data_all[458]);
module_output_bit_459	m459	(input_data_all[1796:0],output_data_all[459]);
module_output_bit_460	m460	(input_data_all[1796:0],output_data_all[460]);
module_output_bit_461	m461	(input_data_all[1796:0],output_data_all[461]);
module_output_bit_462	m462	(input_data_all[1796:0],output_data_all[462]);
module_output_bit_463	m463	(input_data_all[1796:0],output_data_all[463]);
module_output_bit_464	m464	(input_data_all[1796:0],output_data_all[464]);
module_output_bit_465	m465	(input_data_all[1796:0],output_data_all[465]);
module_output_bit_466	m466	(input_data_all[1796:0],output_data_all[466]);
module_output_bit_467	m467	(input_data_all[1796:0],output_data_all[467]);
module_output_bit_468	m468	(input_data_all[1796:0],output_data_all[468]);
module_output_bit_469	m469	(input_data_all[1796:0],output_data_all[469]);
module_output_bit_470	m470	(input_data_all[1796:0],output_data_all[470]);
module_output_bit_471	m471	(input_data_all[1796:0],output_data_all[471]);
module_output_bit_472	m472	(input_data_all[1796:0],output_data_all[472]);
module_output_bit_473	m473	(input_data_all[1796:0],output_data_all[473]);
module_output_bit_474	m474	(input_data_all[1796:0],output_data_all[474]);
module_output_bit_475	m475	(input_data_all[1796:0],output_data_all[475]);
module_output_bit_476	m476	(input_data_all[1796:0],output_data_all[476]);
module_output_bit_477	m477	(input_data_all[1796:0],output_data_all[477]);
module_output_bit_478	m478	(input_data_all[1796:0],output_data_all[478]);
module_output_bit_479	m479	(input_data_all[1796:0],output_data_all[479]);
module_output_bit_480	m480	(input_data_all[1796:0],output_data_all[480]);
module_output_bit_481	m481	(input_data_all[1796:0],output_data_all[481]);
module_output_bit_482	m482	(input_data_all[1796:0],output_data_all[482]);
module_output_bit_483	m483	(input_data_all[1796:0],output_data_all[483]);
module_output_bit_484	m484	(input_data_all[1796:0],output_data_all[484]);
module_output_bit_485	m485	(input_data_all[1796:0],output_data_all[485]);
module_output_bit_486	m486	(input_data_all[1796:0],output_data_all[486]);
module_output_bit_487	m487	(input_data_all[1796:0],output_data_all[487]);
module_output_bit_488	m488	(input_data_all[1796:0],output_data_all[488]);
module_output_bit_489	m489	(input_data_all[1796:0],output_data_all[489]);
module_output_bit_490	m490	(input_data_all[1796:0],output_data_all[490]);
module_output_bit_491	m491	(input_data_all[1796:0],output_data_all[491]);
module_output_bit_492	m492	(input_data_all[1796:0],output_data_all[492]);
module_output_bit_493	m493	(input_data_all[1796:0],output_data_all[493]);
module_output_bit_494	m494	(input_data_all[1796:0],output_data_all[494]);
module_output_bit_495	m495	(input_data_all[1796:0],output_data_all[495]);
module_output_bit_496	m496	(input_data_all[1796:0],output_data_all[496]);
module_output_bit_497	m497	(input_data_all[1796:0],output_data_all[497]);
module_output_bit_498	m498	(input_data_all[1796:0],output_data_all[498]);
module_output_bit_499	m499	(input_data_all[1796:0],output_data_all[499]);
module_output_bit_500	m500	(input_data_all[1796:0],output_data_all[500]);
module_output_bit_501	m501	(input_data_all[1796:0],output_data_all[501]);
module_output_bit_502	m502	(input_data_all[1796:0],output_data_all[502]);
module_output_bit_503	m503	(input_data_all[1796:0],output_data_all[503]);
module_output_bit_504	m504	(input_data_all[1796:0],output_data_all[504]);
module_output_bit_505	m505	(input_data_all[1796:0],output_data_all[505]);
module_output_bit_506	m506	(input_data_all[1796:0],output_data_all[506]);
module_output_bit_507	m507	(input_data_all[1796:0],output_data_all[507]);
module_output_bit_508	m508	(input_data_all[1796:0],output_data_all[508]);
module_output_bit_509	m509	(input_data_all[1796:0],output_data_all[509]);
module_output_bit_510	m510	(input_data_all[1796:0],output_data_all[510]);
module_output_bit_511	m511	(input_data_all[1796:0],output_data_all[511]);
module_output_bit_512	m512	(input_data_all[1796:0],output_data_all[512]);
module_output_bit_513	m513	(input_data_all[1796:0],output_data_all[513]);
module_output_bit_514	m514	(input_data_all[1796:0],output_data_all[514]);
module_output_bit_515	m515	(input_data_all[1796:0],output_data_all[515]);
module_output_bit_516	m516	(input_data_all[1796:0],output_data_all[516]);
module_output_bit_517	m517	(input_data_all[1796:0],output_data_all[517]);
module_output_bit_518	m518	(input_data_all[1796:0],output_data_all[518]);
module_output_bit_519	m519	(input_data_all[1796:0],output_data_all[519]);
module_output_bit_520	m520	(input_data_all[1796:0],output_data_all[520]);
module_output_bit_521	m521	(input_data_all[1796:0],output_data_all[521]);
module_output_bit_522	m522	(input_data_all[1796:0],output_data_all[522]);
module_output_bit_523	m523	(input_data_all[1796:0],output_data_all[523]);
module_output_bit_524	m524	(input_data_all[1796:0],output_data_all[524]);
module_output_bit_525	m525	(input_data_all[1796:0],output_data_all[525]);
module_output_bit_526	m526	(input_data_all[1796:0],output_data_all[526]);
module_output_bit_527	m527	(input_data_all[1796:0],output_data_all[527]);
module_output_bit_528	m528	(input_data_all[1796:0],output_data_all[528]);
module_output_bit_529	m529	(input_data_all[1796:0],output_data_all[529]);
module_output_bit_530	m530	(input_data_all[1796:0],output_data_all[530]);
module_output_bit_531	m531	(input_data_all[1796:0],output_data_all[531]);
module_output_bit_532	m532	(input_data_all[1796:0],output_data_all[532]);
module_output_bit_533	m533	(input_data_all[1796:0],output_data_all[533]);
module_output_bit_534	m534	(input_data_all[1796:0],output_data_all[534]);
module_output_bit_535	m535	(input_data_all[1796:0],output_data_all[535]);
module_output_bit_536	m536	(input_data_all[1796:0],output_data_all[536]);
module_output_bit_537	m537	(input_data_all[1796:0],output_data_all[537]);
module_output_bit_538	m538	(input_data_all[1796:0],output_data_all[538]);
module_output_bit_539	m539	(input_data_all[1796:0],output_data_all[539]);
module_output_bit_540	m540	(input_data_all[1796:0],output_data_all[540]);
module_output_bit_541	m541	(input_data_all[1796:0],output_data_all[541]);
module_output_bit_542	m542	(input_data_all[1796:0],output_data_all[542]);
module_output_bit_543	m543	(input_data_all[1796:0],output_data_all[543]);
module_output_bit_544	m544	(input_data_all[1796:0],output_data_all[544]);
module_output_bit_545	m545	(input_data_all[1796:0],output_data_all[545]);
module_output_bit_546	m546	(input_data_all[1796:0],output_data_all[546]);
module_output_bit_547	m547	(input_data_all[1796:0],output_data_all[547]);
module_output_bit_548	m548	(input_data_all[1796:0],output_data_all[548]);
module_output_bit_549	m549	(input_data_all[1796:0],output_data_all[549]);
module_output_bit_550	m550	(input_data_all[1796:0],output_data_all[550]);
module_output_bit_551	m551	(input_data_all[1796:0],output_data_all[551]);
module_output_bit_552	m552	(input_data_all[1796:0],output_data_all[552]);
module_output_bit_553	m553	(input_data_all[1796:0],output_data_all[553]);
module_output_bit_554	m554	(input_data_all[1796:0],output_data_all[554]);
module_output_bit_555	m555	(input_data_all[1796:0],output_data_all[555]);
module_output_bit_556	m556	(input_data_all[1796:0],output_data_all[556]);
module_output_bit_557	m557	(input_data_all[1796:0],output_data_all[557]);
module_output_bit_558	m558	(input_data_all[1796:0],output_data_all[558]);
module_output_bit_559	m559	(input_data_all[1796:0],output_data_all[559]);
module_output_bit_560	m560	(input_data_all[1796:0],output_data_all[560]);
module_output_bit_561	m561	(input_data_all[1796:0],output_data_all[561]);
module_output_bit_562	m562	(input_data_all[1796:0],output_data_all[562]);
module_output_bit_563	m563	(input_data_all[1796:0],output_data_all[563]);
module_output_bit_564	m564	(input_data_all[1796:0],output_data_all[564]);
module_output_bit_565	m565	(input_data_all[1796:0],output_data_all[565]);
module_output_bit_566	m566	(input_data_all[1796:0],output_data_all[566]);
module_output_bit_567	m567	(input_data_all[1796:0],output_data_all[567]);
module_output_bit_568	m568	(input_data_all[1796:0],output_data_all[568]);
module_output_bit_569	m569	(input_data_all[1796:0],output_data_all[569]);
module_output_bit_570	m570	(input_data_all[1796:0],output_data_all[570]);
module_output_bit_571	m571	(input_data_all[1796:0],output_data_all[571]);
module_output_bit_572	m572	(input_data_all[1796:0],output_data_all[572]);
module_output_bit_573	m573	(input_data_all[1796:0],output_data_all[573]);
module_output_bit_574	m574	(input_data_all[1796:0],output_data_all[574]);
module_output_bit_575	m575	(input_data_all[1796:0],output_data_all[575]);
module_output_bit_576	m576	(input_data_all[1796:0],output_data_all[576]);
module_output_bit_577	m577	(input_data_all[1796:0],output_data_all[577]);
module_output_bit_578	m578	(input_data_all[1796:0],output_data_all[578]);
module_output_bit_579	m579	(input_data_all[1796:0],output_data_all[579]);
module_output_bit_580	m580	(input_data_all[1796:0],output_data_all[580]);
module_output_bit_581	m581	(input_data_all[1796:0],output_data_all[581]);
module_output_bit_582	m582	(input_data_all[1796:0],output_data_all[582]);
module_output_bit_583	m583	(input_data_all[1796:0],output_data_all[583]);
module_output_bit_584	m584	(input_data_all[1796:0],output_data_all[584]);
module_output_bit_585	m585	(input_data_all[1796:0],output_data_all[585]);
module_output_bit_586	m586	(input_data_all[1796:0],output_data_all[586]);
module_output_bit_587	m587	(input_data_all[1796:0],output_data_all[587]);
module_output_bit_588	m588	(input_data_all[1796:0],output_data_all[588]);
module_output_bit_589	m589	(input_data_all[1796:0],output_data_all[589]);
module_output_bit_590	m590	(input_data_all[1796:0],output_data_all[590]);
module_output_bit_591	m591	(input_data_all[1796:0],output_data_all[591]);
module_output_bit_592	m592	(input_data_all[1796:0],output_data_all[592]);
module_output_bit_593	m593	(input_data_all[1796:0],output_data_all[593]);
module_output_bit_594	m594	(input_data_all[1796:0],output_data_all[594]);
module_output_bit_595	m595	(input_data_all[1796:0],output_data_all[595]);
module_output_bit_596	m596	(input_data_all[1796:0],output_data_all[596]);
module_output_bit_597	m597	(input_data_all[1796:0],output_data_all[597]);
module_output_bit_598	m598	(input_data_all[1796:0],output_data_all[598]);
module_output_bit_599	m599	(input_data_all[1796:0],output_data_all[599]);
module_output_bit_600	m600	(input_data_all[1796:0],output_data_all[600]);
module_output_bit_601	m601	(input_data_all[1796:0],output_data_all[601]);
module_output_bit_602	m602	(input_data_all[1796:0],output_data_all[602]);
module_output_bit_603	m603	(input_data_all[1796:0],output_data_all[603]);
module_output_bit_604	m604	(input_data_all[1796:0],output_data_all[604]);
module_output_bit_605	m605	(input_data_all[1796:0],output_data_all[605]);
module_output_bit_606	m606	(input_data_all[1796:0],output_data_all[606]);
module_output_bit_607	m607	(input_data_all[1796:0],output_data_all[607]);
module_output_bit_608	m608	(input_data_all[1796:0],output_data_all[608]);
module_output_bit_609	m609	(input_data_all[1796:0],output_data_all[609]);
module_output_bit_610	m610	(input_data_all[1796:0],output_data_all[610]);
module_output_bit_611	m611	(input_data_all[1796:0],output_data_all[611]);
module_output_bit_612	m612	(input_data_all[1796:0],output_data_all[612]);
module_output_bit_613	m613	(input_data_all[1796:0],output_data_all[613]);
module_output_bit_614	m614	(input_data_all[1796:0],output_data_all[614]);
module_output_bit_615	m615	(input_data_all[1796:0],output_data_all[615]);
module_output_bit_616	m616	(input_data_all[1796:0],output_data_all[616]);
module_output_bit_617	m617	(input_data_all[1796:0],output_data_all[617]);
module_output_bit_618	m618	(input_data_all[1796:0],output_data_all[618]);
module_output_bit_619	m619	(input_data_all[1796:0],output_data_all[619]);
module_output_bit_620	m620	(input_data_all[1796:0],output_data_all[620]);
module_output_bit_621	m621	(input_data_all[1796:0],output_data_all[621]);
module_output_bit_622	m622	(input_data_all[1796:0],output_data_all[622]);
module_output_bit_623	m623	(input_data_all[1796:0],output_data_all[623]);
module_output_bit_624	m624	(input_data_all[1796:0],output_data_all[624]);
module_output_bit_625	m625	(input_data_all[1796:0],output_data_all[625]);
module_output_bit_626	m626	(input_data_all[1796:0],output_data_all[626]);
module_output_bit_627	m627	(input_data_all[1796:0],output_data_all[627]);
module_output_bit_628	m628	(input_data_all[1796:0],output_data_all[628]);
module_output_bit_629	m629	(input_data_all[1796:0],output_data_all[629]);
module_output_bit_630	m630	(input_data_all[1796:0],output_data_all[630]);
module_output_bit_631	m631	(input_data_all[1796:0],output_data_all[631]);
module_output_bit_632	m632	(input_data_all[1796:0],output_data_all[632]);
module_output_bit_633	m633	(input_data_all[1796:0],output_data_all[633]);
module_output_bit_634	m634	(input_data_all[1796:0],output_data_all[634]);
module_output_bit_635	m635	(input_data_all[1796:0],output_data_all[635]);
module_output_bit_636	m636	(input_data_all[1796:0],output_data_all[636]);
module_output_bit_637	m637	(input_data_all[1796:0],output_data_all[637]);
module_output_bit_638	m638	(input_data_all[1796:0],output_data_all[638]);
module_output_bit_639	m639	(input_data_all[1796:0],output_data_all[639]);
module_output_bit_640	m640	(input_data_all[1796:0],output_data_all[640]);
module_output_bit_641	m641	(input_data_all[1796:0],output_data_all[641]);
module_output_bit_642	m642	(input_data_all[1796:0],output_data_all[642]);
module_output_bit_643	m643	(input_data_all[1796:0],output_data_all[643]);
module_output_bit_644	m644	(input_data_all[1796:0],output_data_all[644]);
module_output_bit_645	m645	(input_data_all[1796:0],output_data_all[645]);
module_output_bit_646	m646	(input_data_all[1796:0],output_data_all[646]);
module_output_bit_647	m647	(input_data_all[1796:0],output_data_all[647]);
module_output_bit_648	m648	(input_data_all[1796:0],output_data_all[648]);
module_output_bit_649	m649	(input_data_all[1796:0],output_data_all[649]);
module_output_bit_650	m650	(input_data_all[1796:0],output_data_all[650]);
module_output_bit_651	m651	(input_data_all[1796:0],output_data_all[651]);
module_output_bit_652	m652	(input_data_all[1796:0],output_data_all[652]);
module_output_bit_653	m653	(input_data_all[1796:0],output_data_all[653]);
module_output_bit_654	m654	(input_data_all[1796:0],output_data_all[654]);
module_output_bit_655	m655	(input_data_all[1796:0],output_data_all[655]);
module_output_bit_656	m656	(input_data_all[1796:0],output_data_all[656]);
module_output_bit_657	m657	(input_data_all[1796:0],output_data_all[657]);
module_output_bit_658	m658	(input_data_all[1796:0],output_data_all[658]);
module_output_bit_659	m659	(input_data_all[1796:0],output_data_all[659]);
module_output_bit_660	m660	(input_data_all[1796:0],output_data_all[660]);
module_output_bit_661	m661	(input_data_all[1796:0],output_data_all[661]);
module_output_bit_662	m662	(input_data_all[1796:0],output_data_all[662]);
module_output_bit_663	m663	(input_data_all[1796:0],output_data_all[663]);
module_output_bit_664	m664	(input_data_all[1796:0],output_data_all[664]);
module_output_bit_665	m665	(input_data_all[1796:0],output_data_all[665]);
module_output_bit_666	m666	(input_data_all[1796:0],output_data_all[666]);
module_output_bit_667	m667	(input_data_all[1796:0],output_data_all[667]);
module_output_bit_668	m668	(input_data_all[1796:0],output_data_all[668]);
module_output_bit_669	m669	(input_data_all[1796:0],output_data_all[669]);
module_output_bit_670	m670	(input_data_all[1796:0],output_data_all[670]);
module_output_bit_671	m671	(input_data_all[1796:0],output_data_all[671]);
module_output_bit_672	m672	(input_data_all[1796:0],output_data_all[672]);
module_output_bit_673	m673	(input_data_all[1796:0],output_data_all[673]);
module_output_bit_674	m674	(input_data_all[1796:0],output_data_all[674]);
module_output_bit_675	m675	(input_data_all[1796:0],output_data_all[675]);
module_output_bit_676	m676	(input_data_all[1796:0],output_data_all[676]);
module_output_bit_677	m677	(input_data_all[1796:0],output_data_all[677]);
module_output_bit_678	m678	(input_data_all[1796:0],output_data_all[678]);
module_output_bit_679	m679	(input_data_all[1796:0],output_data_all[679]);
module_output_bit_680	m680	(input_data_all[1796:0],output_data_all[680]);
module_output_bit_681	m681	(input_data_all[1796:0],output_data_all[681]);
module_output_bit_682	m682	(input_data_all[1796:0],output_data_all[682]);
module_output_bit_683	m683	(input_data_all[1796:0],output_data_all[683]);
module_output_bit_684	m684	(input_data_all[1796:0],output_data_all[684]);
module_output_bit_685	m685	(input_data_all[1796:0],output_data_all[685]);
module_output_bit_686	m686	(input_data_all[1796:0],output_data_all[686]);
module_output_bit_687	m687	(input_data_all[1796:0],output_data_all[687]);
module_output_bit_688	m688	(input_data_all[1796:0],output_data_all[688]);
module_output_bit_689	m689	(input_data_all[1796:0],output_data_all[689]);
module_output_bit_690	m690	(input_data_all[1796:0],output_data_all[690]);
module_output_bit_691	m691	(input_data_all[1796:0],output_data_all[691]);
module_output_bit_692	m692	(input_data_all[1796:0],output_data_all[692]);
module_output_bit_693	m693	(input_data_all[1796:0],output_data_all[693]);
module_output_bit_694	m694	(input_data_all[1796:0],output_data_all[694]);
module_output_bit_695	m695	(input_data_all[1796:0],output_data_all[695]);
module_output_bit_696	m696	(input_data_all[1796:0],output_data_all[696]);
module_output_bit_697	m697	(input_data_all[1796:0],output_data_all[697]);
module_output_bit_698	m698	(input_data_all[1796:0],output_data_all[698]);
module_output_bit_699	m699	(input_data_all[1796:0],output_data_all[699]);
module_output_bit_700	m700	(input_data_all[1796:0],output_data_all[700]);
module_output_bit_701	m701	(input_data_all[1796:0],output_data_all[701]);
module_output_bit_702	m702	(input_data_all[1796:0],output_data_all[702]);
module_output_bit_703	m703	(input_data_all[1796:0],output_data_all[703]);
module_output_bit_704	m704	(input_data_all[1796:0],output_data_all[704]);
module_output_bit_705	m705	(input_data_all[1796:0],output_data_all[705]);
module_output_bit_706	m706	(input_data_all[1796:0],output_data_all[706]);
module_output_bit_707	m707	(input_data_all[1796:0],output_data_all[707]);
module_output_bit_708	m708	(input_data_all[1796:0],output_data_all[708]);
module_output_bit_709	m709	(input_data_all[1796:0],output_data_all[709]);
module_output_bit_710	m710	(input_data_all[1796:0],output_data_all[710]);
module_output_bit_711	m711	(input_data_all[1796:0],output_data_all[711]);
module_output_bit_712	m712	(input_data_all[1796:0],output_data_all[712]);
module_output_bit_713	m713	(input_data_all[1796:0],output_data_all[713]);
module_output_bit_714	m714	(input_data_all[1796:0],output_data_all[714]);
module_output_bit_715	m715	(input_data_all[1796:0],output_data_all[715]);
module_output_bit_716	m716	(input_data_all[1796:0],output_data_all[716]);
module_output_bit_717	m717	(input_data_all[1796:0],output_data_all[717]);
module_output_bit_718	m718	(input_data_all[1796:0],output_data_all[718]);
module_output_bit_719	m719	(input_data_all[1796:0],output_data_all[719]);
module_output_bit_720	m720	(input_data_all[1796:0],output_data_all[720]);
module_output_bit_721	m721	(input_data_all[1796:0],output_data_all[721]);
module_output_bit_722	m722	(input_data_all[1796:0],output_data_all[722]);
module_output_bit_723	m723	(input_data_all[1796:0],output_data_all[723]);
module_output_bit_724	m724	(input_data_all[1796:0],output_data_all[724]);
module_output_bit_725	m725	(input_data_all[1796:0],output_data_all[725]);
module_output_bit_726	m726	(input_data_all[1796:0],output_data_all[726]);
module_output_bit_727	m727	(input_data_all[1796:0],output_data_all[727]);
module_output_bit_728	m728	(input_data_all[1796:0],output_data_all[728]);
module_output_bit_729	m729	(input_data_all[1796:0],output_data_all[729]);
module_output_bit_730	m730	(input_data_all[1796:0],output_data_all[730]);
module_output_bit_731	m731	(input_data_all[1796:0],output_data_all[731]);
module_output_bit_732	m732	(input_data_all[1796:0],output_data_all[732]);
module_output_bit_733	m733	(input_data_all[1796:0],output_data_all[733]);
module_output_bit_734	m734	(input_data_all[1796:0],output_data_all[734]);
module_output_bit_735	m735	(input_data_all[1796:0],output_data_all[735]);
module_output_bit_736	m736	(input_data_all[1796:0],output_data_all[736]);
module_output_bit_737	m737	(input_data_all[1796:0],output_data_all[737]);
module_output_bit_738	m738	(input_data_all[1796:0],output_data_all[738]);
module_output_bit_739	m739	(input_data_all[1796:0],output_data_all[739]);
module_output_bit_740	m740	(input_data_all[1796:0],output_data_all[740]);
module_output_bit_741	m741	(input_data_all[1796:0],output_data_all[741]);
module_output_bit_742	m742	(input_data_all[1796:0],output_data_all[742]);
module_output_bit_743	m743	(input_data_all[1796:0],output_data_all[743]);
module_output_bit_744	m744	(input_data_all[1796:0],output_data_all[744]);
module_output_bit_745	m745	(input_data_all[1796:0],output_data_all[745]);
module_output_bit_746	m746	(input_data_all[1796:0],output_data_all[746]);
module_output_bit_747	m747	(input_data_all[1796:0],output_data_all[747]);
module_output_bit_748	m748	(input_data_all[1796:0],output_data_all[748]);
module_output_bit_749	m749	(input_data_all[1796:0],output_data_all[749]);
module_output_bit_750	m750	(input_data_all[1796:0],output_data_all[750]);
module_output_bit_751	m751	(input_data_all[1796:0],output_data_all[751]);
module_output_bit_752	m752	(input_data_all[1796:0],output_data_all[752]);
module_output_bit_753	m753	(input_data_all[1796:0],output_data_all[753]);
module_output_bit_754	m754	(input_data_all[1796:0],output_data_all[754]);
module_output_bit_755	m755	(input_data_all[1796:0],output_data_all[755]);
module_output_bit_756	m756	(input_data_all[1796:0],output_data_all[756]);
module_output_bit_757	m757	(input_data_all[1796:0],output_data_all[757]);
module_output_bit_758	m758	(input_data_all[1796:0],output_data_all[758]);
module_output_bit_759	m759	(input_data_all[1796:0],output_data_all[759]);
module_output_bit_760	m760	(input_data_all[1796:0],output_data_all[760]);
module_output_bit_761	m761	(input_data_all[1796:0],output_data_all[761]);
module_output_bit_762	m762	(input_data_all[1796:0],output_data_all[762]);
module_output_bit_763	m763	(input_data_all[1796:0],output_data_all[763]);
module_output_bit_764	m764	(input_data_all[1796:0],output_data_all[764]);
module_output_bit_765	m765	(input_data_all[1796:0],output_data_all[765]);
module_output_bit_766	m766	(input_data_all[1796:0],output_data_all[766]);
module_output_bit_767	m767	(input_data_all[1796:0],output_data_all[767]);
module_output_bit_768	m768	(input_data_all[1796:0],output_data_all[768]);
module_output_bit_769	m769	(input_data_all[1796:0],output_data_all[769]);
module_output_bit_770	m770	(input_data_all[1796:0],output_data_all[770]);
module_output_bit_771	m771	(input_data_all[1796:0],output_data_all[771]);
module_output_bit_772	m772	(input_data_all[1796:0],output_data_all[772]);
module_output_bit_773	m773	(input_data_all[1796:0],output_data_all[773]);
module_output_bit_774	m774	(input_data_all[1796:0],output_data_all[774]);
module_output_bit_775	m775	(input_data_all[1796:0],output_data_all[775]);
module_output_bit_776	m776	(input_data_all[1796:0],output_data_all[776]);
module_output_bit_777	m777	(input_data_all[1796:0],output_data_all[777]);
module_output_bit_778	m778	(input_data_all[1796:0],output_data_all[778]);
module_output_bit_779	m779	(input_data_all[1796:0],output_data_all[779]);
module_output_bit_780	m780	(input_data_all[1796:0],output_data_all[780]);
module_output_bit_781	m781	(input_data_all[1796:0],output_data_all[781]);
module_output_bit_782	m782	(input_data_all[1796:0],output_data_all[782]);
module_output_bit_783	m783	(input_data_all[1796:0],output_data_all[783]);
module_output_bit_784	m784	(input_data_all[1796:0],output_data_all[784]);
module_output_bit_785	m785	(input_data_all[1796:0],output_data_all[785]);
module_output_bit_786	m786	(input_data_all[1796:0],output_data_all[786]);
module_output_bit_787	m787	(input_data_all[1796:0],output_data_all[787]);
module_output_bit_788	m788	(input_data_all[1796:0],output_data_all[788]);
module_output_bit_789	m789	(input_data_all[1796:0],output_data_all[789]);
module_output_bit_790	m790	(input_data_all[1796:0],output_data_all[790]);
module_output_bit_791	m791	(input_data_all[1796:0],output_data_all[791]);
module_output_bit_792	m792	(input_data_all[1796:0],output_data_all[792]);
module_output_bit_793	m793	(input_data_all[1796:0],output_data_all[793]);
module_output_bit_794	m794	(input_data_all[1796:0],output_data_all[794]);
module_output_bit_795	m795	(input_data_all[1796:0],output_data_all[795]);
module_output_bit_796	m796	(input_data_all[1796:0],output_data_all[796]);
module_output_bit_797	m797	(input_data_all[1796:0],output_data_all[797]);
module_output_bit_798	m798	(input_data_all[1796:0],output_data_all[798]);
module_output_bit_799	m799	(input_data_all[1796:0],output_data_all[799]);
module_output_bit_800	m800	(input_data_all[1796:0],output_data_all[800]);
module_output_bit_801	m801	(input_data_all[1796:0],output_data_all[801]);
module_output_bit_802	m802	(input_data_all[1796:0],output_data_all[802]);
module_output_bit_803	m803	(input_data_all[1796:0],output_data_all[803]);
module_output_bit_804	m804	(input_data_all[1796:0],output_data_all[804]);
module_output_bit_805	m805	(input_data_all[1796:0],output_data_all[805]);
module_output_bit_806	m806	(input_data_all[1796:0],output_data_all[806]);
module_output_bit_807	m807	(input_data_all[1796:0],output_data_all[807]);
module_output_bit_808	m808	(input_data_all[1796:0],output_data_all[808]);
module_output_bit_809	m809	(input_data_all[1796:0],output_data_all[809]);
module_output_bit_810	m810	(input_data_all[1796:0],output_data_all[810]);
module_output_bit_811	m811	(input_data_all[1796:0],output_data_all[811]);
module_output_bit_812	m812	(input_data_all[1796:0],output_data_all[812]);
module_output_bit_813	m813	(input_data_all[1796:0],output_data_all[813]);
module_output_bit_814	m814	(input_data_all[1796:0],output_data_all[814]);
module_output_bit_815	m815	(input_data_all[1796:0],output_data_all[815]);
module_output_bit_816	m816	(input_data_all[1796:0],output_data_all[816]);
module_output_bit_817	m817	(input_data_all[1796:0],output_data_all[817]);
module_output_bit_818	m818	(input_data_all[1796:0],output_data_all[818]);
module_output_bit_819	m819	(input_data_all[1796:0],output_data_all[819]);
module_output_bit_820	m820	(input_data_all[1796:0],output_data_all[820]);
module_output_bit_821	m821	(input_data_all[1796:0],output_data_all[821]);
module_output_bit_822	m822	(input_data_all[1796:0],output_data_all[822]);
module_output_bit_823	m823	(input_data_all[1796:0],output_data_all[823]);
module_output_bit_824	m824	(input_data_all[1796:0],output_data_all[824]);
module_output_bit_825	m825	(input_data_all[1796:0],output_data_all[825]);
module_output_bit_826	m826	(input_data_all[1796:0],output_data_all[826]);
module_output_bit_827	m827	(input_data_all[1796:0],output_data_all[827]);
module_output_bit_828	m828	(input_data_all[1796:0],output_data_all[828]);
module_output_bit_829	m829	(input_data_all[1796:0],output_data_all[829]);
module_output_bit_830	m830	(input_data_all[1796:0],output_data_all[830]);
module_output_bit_831	m831	(input_data_all[1796:0],output_data_all[831]);
module_output_bit_832	m832	(input_data_all[1796:0],output_data_all[832]);
module_output_bit_833	m833	(input_data_all[1796:0],output_data_all[833]);
module_output_bit_834	m834	(input_data_all[1796:0],output_data_all[834]);
module_output_bit_835	m835	(input_data_all[1796:0],output_data_all[835]);
module_output_bit_836	m836	(input_data_all[1796:0],output_data_all[836]);
module_output_bit_837	m837	(input_data_all[1796:0],output_data_all[837]);
module_output_bit_838	m838	(input_data_all[1796:0],output_data_all[838]);
module_output_bit_839	m839	(input_data_all[1796:0],output_data_all[839]);
module_output_bit_840	m840	(input_data_all[1796:0],output_data_all[840]);
module_output_bit_841	m841	(input_data_all[1796:0],output_data_all[841]);
module_output_bit_842	m842	(input_data_all[1796:0],output_data_all[842]);
module_output_bit_843	m843	(input_data_all[1796:0],output_data_all[843]);
module_output_bit_844	m844	(input_data_all[1796:0],output_data_all[844]);
module_output_bit_845	m845	(input_data_all[1796:0],output_data_all[845]);
module_output_bit_846	m846	(input_data_all[1796:0],output_data_all[846]);
module_output_bit_847	m847	(input_data_all[1796:0],output_data_all[847]);
module_output_bit_848	m848	(input_data_all[1796:0],output_data_all[848]);
module_output_bit_849	m849	(input_data_all[1796:0],output_data_all[849]);
module_output_bit_850	m850	(input_data_all[1796:0],output_data_all[850]);
module_output_bit_851	m851	(input_data_all[1796:0],output_data_all[851]);
module_output_bit_852	m852	(input_data_all[1796:0],output_data_all[852]);
module_output_bit_853	m853	(input_data_all[1796:0],output_data_all[853]);
module_output_bit_854	m854	(input_data_all[1796:0],output_data_all[854]);
module_output_bit_855	m855	(input_data_all[1796:0],output_data_all[855]);
module_output_bit_856	m856	(input_data_all[1796:0],output_data_all[856]);
module_output_bit_857	m857	(input_data_all[1796:0],output_data_all[857]);
module_output_bit_858	m858	(input_data_all[1796:0],output_data_all[858]);
module_output_bit_859	m859	(input_data_all[1796:0],output_data_all[859]);
module_output_bit_860	m860	(input_data_all[1796:0],output_data_all[860]);
module_output_bit_861	m861	(input_data_all[1796:0],output_data_all[861]);
module_output_bit_862	m862	(input_data_all[1796:0],output_data_all[862]);
module_output_bit_863	m863	(input_data_all[1796:0],output_data_all[863]);
module_output_bit_864	m864	(input_data_all[1796:0],output_data_all[864]);
module_output_bit_865	m865	(input_data_all[1796:0],output_data_all[865]);
module_output_bit_866	m866	(input_data_all[1796:0],output_data_all[866]);
module_output_bit_867	m867	(input_data_all[1796:0],output_data_all[867]);
module_output_bit_868	m868	(input_data_all[1796:0],output_data_all[868]);
module_output_bit_869	m869	(input_data_all[1796:0],output_data_all[869]);
module_output_bit_870	m870	(input_data_all[1796:0],output_data_all[870]);
module_output_bit_871	m871	(input_data_all[1796:0],output_data_all[871]);
module_output_bit_872	m872	(input_data_all[1796:0],output_data_all[872]);
module_output_bit_873	m873	(input_data_all[1796:0],output_data_all[873]);
module_output_bit_874	m874	(input_data_all[1796:0],output_data_all[874]);
module_output_bit_875	m875	(input_data_all[1796:0],output_data_all[875]);
module_output_bit_876	m876	(input_data_all[1796:0],output_data_all[876]);
module_output_bit_877	m877	(input_data_all[1796:0],output_data_all[877]);
module_output_bit_878	m878	(input_data_all[1796:0],output_data_all[878]);
module_output_bit_879	m879	(input_data_all[1796:0],output_data_all[879]);
module_output_bit_880	m880	(input_data_all[1796:0],output_data_all[880]);
module_output_bit_881	m881	(input_data_all[1796:0],output_data_all[881]);
module_output_bit_882	m882	(input_data_all[1796:0],output_data_all[882]);
module_output_bit_883	m883	(input_data_all[1796:0],output_data_all[883]);
module_output_bit_884	m884	(input_data_all[1796:0],output_data_all[884]);
module_output_bit_885	m885	(input_data_all[1796:0],output_data_all[885]);
module_output_bit_886	m886	(input_data_all[1796:0],output_data_all[886]);
module_output_bit_887	m887	(input_data_all[1796:0],output_data_all[887]);
module_output_bit_888	m888	(input_data_all[1796:0],output_data_all[888]);
module_output_bit_889	m889	(input_data_all[1796:0],output_data_all[889]);
module_output_bit_890	m890	(input_data_all[1796:0],output_data_all[890]);
module_output_bit_891	m891	(input_data_all[1796:0],output_data_all[891]);
module_output_bit_892	m892	(input_data_all[1796:0],output_data_all[892]);
module_output_bit_893	m893	(input_data_all[1796:0],output_data_all[893]);
module_output_bit_894	m894	(input_data_all[1796:0],output_data_all[894]);
module_output_bit_895	m895	(input_data_all[1796:0],output_data_all[895]);
module_output_bit_896	m896	(input_data_all[1796:0],output_data_all[896]);
module_output_bit_897	m897	(input_data_all[1796:0],output_data_all[897]);
module_output_bit_898	m898	(input_data_all[1796:0],output_data_all[898]);
module_output_bit_899	m899	(input_data_all[1796:0],output_data_all[899]);
module_output_bit_900	m900	(input_data_all[1796:0],output_data_all[900]);
module_output_bit_901	m901	(input_data_all[1796:0],output_data_all[901]);
module_output_bit_902	m902	(input_data_all[1796:0],output_data_all[902]);
module_output_bit_903	m903	(input_data_all[1796:0],output_data_all[903]);
module_output_bit_904	m904	(input_data_all[1796:0],output_data_all[904]);
module_output_bit_905	m905	(input_data_all[1796:0],output_data_all[905]);
module_output_bit_906	m906	(input_data_all[1796:0],output_data_all[906]);
module_output_bit_907	m907	(input_data_all[1796:0],output_data_all[907]);
module_output_bit_908	m908	(input_data_all[1796:0],output_data_all[908]);
module_output_bit_909	m909	(input_data_all[1796:0],output_data_all[909]);
module_output_bit_910	m910	(input_data_all[1796:0],output_data_all[910]);
module_output_bit_911	m911	(input_data_all[1796:0],output_data_all[911]);
module_output_bit_912	m912	(input_data_all[1796:0],output_data_all[912]);
module_output_bit_913	m913	(input_data_all[1796:0],output_data_all[913]);
module_output_bit_914	m914	(input_data_all[1796:0],output_data_all[914]);
module_output_bit_915	m915	(input_data_all[1796:0],output_data_all[915]);
module_output_bit_916	m916	(input_data_all[1796:0],output_data_all[916]);
module_output_bit_917	m917	(input_data_all[1796:0],output_data_all[917]);
module_output_bit_918	m918	(input_data_all[1796:0],output_data_all[918]);
module_output_bit_919	m919	(input_data_all[1796:0],output_data_all[919]);
module_output_bit_920	m920	(input_data_all[1796:0],output_data_all[920]);
module_output_bit_921	m921	(input_data_all[1796:0],output_data_all[921]);
module_output_bit_922	m922	(input_data_all[1796:0],output_data_all[922]);
module_output_bit_923	m923	(input_data_all[1796:0],output_data_all[923]);
module_output_bit_924	m924	(input_data_all[1796:0],output_data_all[924]);
module_output_bit_925	m925	(input_data_all[1796:0],output_data_all[925]);
module_output_bit_926	m926	(input_data_all[1796:0],output_data_all[926]);
module_output_bit_927	m927	(input_data_all[1796:0],output_data_all[927]);
module_output_bit_928	m928	(input_data_all[1796:0],output_data_all[928]);
module_output_bit_929	m929	(input_data_all[1796:0],output_data_all[929]);
module_output_bit_930	m930	(input_data_all[1796:0],output_data_all[930]);
module_output_bit_931	m931	(input_data_all[1796:0],output_data_all[931]);
module_output_bit_932	m932	(input_data_all[1796:0],output_data_all[932]);
module_output_bit_933	m933	(input_data_all[1796:0],output_data_all[933]);
module_output_bit_934	m934	(input_data_all[1796:0],output_data_all[934]);
module_output_bit_935	m935	(input_data_all[1796:0],output_data_all[935]);
module_output_bit_936	m936	(input_data_all[1796:0],output_data_all[936]);
module_output_bit_937	m937	(input_data_all[1796:0],output_data_all[937]);
module_output_bit_938	m938	(input_data_all[1796:0],output_data_all[938]);
module_output_bit_939	m939	(input_data_all[1796:0],output_data_all[939]);
module_output_bit_940	m940	(input_data_all[1796:0],output_data_all[940]);
module_output_bit_941	m941	(input_data_all[1796:0],output_data_all[941]);
module_output_bit_942	m942	(input_data_all[1796:0],output_data_all[942]);
module_output_bit_943	m943	(input_data_all[1796:0],output_data_all[943]);
module_output_bit_944	m944	(input_data_all[1796:0],output_data_all[944]);
module_output_bit_945	m945	(input_data_all[1796:0],output_data_all[945]);
module_output_bit_946	m946	(input_data_all[1796:0],output_data_all[946]);
module_output_bit_947	m947	(input_data_all[1796:0],output_data_all[947]);
module_output_bit_948	m948	(input_data_all[1796:0],output_data_all[948]);
module_output_bit_949	m949	(input_data_all[1796:0],output_data_all[949]);
module_output_bit_950	m950	(input_data_all[1796:0],output_data_all[950]);
module_output_bit_951	m951	(input_data_all[1796:0],output_data_all[951]);
module_output_bit_952	m952	(input_data_all[1796:0],output_data_all[952]);
module_output_bit_953	m953	(input_data_all[1796:0],output_data_all[953]);
module_output_bit_954	m954	(input_data_all[1796:0],output_data_all[954]);
module_output_bit_955	m955	(input_data_all[1796:0],output_data_all[955]);
module_output_bit_956	m956	(input_data_all[1796:0],output_data_all[956]);
module_output_bit_957	m957	(input_data_all[1796:0],output_data_all[957]);
module_output_bit_958	m958	(input_data_all[1796:0],output_data_all[958]);
module_output_bit_959	m959	(input_data_all[1796:0],output_data_all[959]);
module_output_bit_960	m960	(input_data_all[1796:0],output_data_all[960]);
module_output_bit_961	m961	(input_data_all[1796:0],output_data_all[961]);
module_output_bit_962	m962	(input_data_all[1796:0],output_data_all[962]);
module_output_bit_963	m963	(input_data_all[1796:0],output_data_all[963]);
module_output_bit_964	m964	(input_data_all[1796:0],output_data_all[964]);
module_output_bit_965	m965	(input_data_all[1796:0],output_data_all[965]);
module_output_bit_966	m966	(input_data_all[1796:0],output_data_all[966]);
module_output_bit_967	m967	(input_data_all[1796:0],output_data_all[967]);
module_output_bit_968	m968	(input_data_all[1796:0],output_data_all[968]);
module_output_bit_969	m969	(input_data_all[1796:0],output_data_all[969]);
module_output_bit_970	m970	(input_data_all[1796:0],output_data_all[970]);
module_output_bit_971	m971	(input_data_all[1796:0],output_data_all[971]);
module_output_bit_972	m972	(input_data_all[1796:0],output_data_all[972]);
module_output_bit_973	m973	(input_data_all[1796:0],output_data_all[973]);
module_output_bit_974	m974	(input_data_all[1796:0],output_data_all[974]);
module_output_bit_975	m975	(input_data_all[1796:0],output_data_all[975]);
module_output_bit_976	m976	(input_data_all[1796:0],output_data_all[976]);
module_output_bit_977	m977	(input_data_all[1796:0],output_data_all[977]);
module_output_bit_978	m978	(input_data_all[1796:0],output_data_all[978]);
module_output_bit_979	m979	(input_data_all[1796:0],output_data_all[979]);
module_output_bit_980	m980	(input_data_all[1796:0],output_data_all[980]);
module_output_bit_981	m981	(input_data_all[1796:0],output_data_all[981]);
module_output_bit_982	m982	(input_data_all[1796:0],output_data_all[982]);
module_output_bit_983	m983	(input_data_all[1796:0],output_data_all[983]);
module_output_bit_984	m984	(input_data_all[1796:0],output_data_all[984]);
module_output_bit_985	m985	(input_data_all[1796:0],output_data_all[985]);
module_output_bit_986	m986	(input_data_all[1796:0],output_data_all[986]);
module_output_bit_987	m987	(input_data_all[1796:0],output_data_all[987]);
module_output_bit_988	m988	(input_data_all[1796:0],output_data_all[988]);
module_output_bit_989	m989	(input_data_all[1796:0],output_data_all[989]);
module_output_bit_990	m990	(input_data_all[1796:0],output_data_all[990]);
module_output_bit_991	m991	(input_data_all[1796:0],output_data_all[991]);
module_output_bit_992	m992	(input_data_all[1796:0],output_data_all[992]);
module_output_bit_993	m993	(input_data_all[1796:0],output_data_all[993]);
module_output_bit_994	m994	(input_data_all[1796:0],output_data_all[994]);
module_output_bit_995	m995	(input_data_all[1796:0],output_data_all[995]);
module_output_bit_996	m996	(input_data_all[1796:0],output_data_all[996]);
module_output_bit_997	m997	(input_data_all[1796:0],output_data_all[997]);
module_output_bit_998	m998	(input_data_all[1796:0],output_data_all[998]);
module_output_bit_999	m999	(input_data_all[1796:0],output_data_all[999]);
module_output_bit_1000	m1000	(input_data_all[1796:0],output_data_all[1000]);
module_output_bit_1001	m1001	(input_data_all[1796:0],output_data_all[1001]);
module_output_bit_1002	m1002	(input_data_all[1796:0],output_data_all[1002]);
module_output_bit_1003	m1003	(input_data_all[1796:0],output_data_all[1003]);
module_output_bit_1004	m1004	(input_data_all[1796:0],output_data_all[1004]);
module_output_bit_1005	m1005	(input_data_all[1796:0],output_data_all[1005]);
module_output_bit_1006	m1006	(input_data_all[1796:0],output_data_all[1006]);
module_output_bit_1007	m1007	(input_data_all[1796:0],output_data_all[1007]);
module_output_bit_1008	m1008	(input_data_all[1796:0],output_data_all[1008]);
module_output_bit_1009	m1009	(input_data_all[1796:0],output_data_all[1009]);
module_output_bit_1010	m1010	(input_data_all[1796:0],output_data_all[1010]);
module_output_bit_1011	m1011	(input_data_all[1796:0],output_data_all[1011]);
module_output_bit_1012	m1012	(input_data_all[1796:0],output_data_all[1012]);
module_output_bit_1013	m1013	(input_data_all[1796:0],output_data_all[1013]);
module_output_bit_1014	m1014	(input_data_all[1796:0],output_data_all[1014]);
module_output_bit_1015	m1015	(input_data_all[1796:0],output_data_all[1015]);
module_output_bit_1016	m1016	(input_data_all[1796:0],output_data_all[1016]);
module_output_bit_1017	m1017	(input_data_all[1796:0],output_data_all[1017]);
module_output_bit_1018	m1018	(input_data_all[1796:0],output_data_all[1018]);
module_output_bit_1019	m1019	(input_data_all[1796:0],output_data_all[1019]);
module_output_bit_1020	m1020	(input_data_all[1796:0],output_data_all[1020]);
module_output_bit_1021	m1021	(input_data_all[1796:0],output_data_all[1021]);
module_output_bit_1022	m1022	(input_data_all[1796:0],output_data_all[1022]);
module_output_bit_1023	m1023	(input_data_all[1796:0],output_data_all[1023]);
module_output_bit_1024	m1024	(input_data_all[1796:0],output_data_all[1024]);
module_output_bit_1025	m1025	(input_data_all[1796:0],output_data_all[1025]);
module_output_bit_1026	m1026	(input_data_all[1796:0],output_data_all[1026]);
module_output_bit_1027	m1027	(input_data_all[1796:0],output_data_all[1027]);
module_output_bit_1028	m1028	(input_data_all[1796:0],output_data_all[1028]);
module_output_bit_1029	m1029	(input_data_all[1796:0],output_data_all[1029]);
module_output_bit_1030	m1030	(input_data_all[1796:0],output_data_all[1030]);
module_output_bit_1031	m1031	(input_data_all[1796:0],output_data_all[1031]);
module_output_bit_1032	m1032	(input_data_all[1796:0],output_data_all[1032]);
module_output_bit_1033	m1033	(input_data_all[1796:0],output_data_all[1033]);
module_output_bit_1034	m1034	(input_data_all[1796:0],output_data_all[1034]);
module_output_bit_1035	m1035	(input_data_all[1796:0],output_data_all[1035]);
module_output_bit_1036	m1036	(input_data_all[1796:0],output_data_all[1036]);
module_output_bit_1037	m1037	(input_data_all[1796:0],output_data_all[1037]);
module_output_bit_1038	m1038	(input_data_all[1796:0],output_data_all[1038]);
module_output_bit_1039	m1039	(input_data_all[1796:0],output_data_all[1039]);
module_output_bit_1040	m1040	(input_data_all[1796:0],output_data_all[1040]);
module_output_bit_1041	m1041	(input_data_all[1796:0],output_data_all[1041]);
module_output_bit_1042	m1042	(input_data_all[1796:0],output_data_all[1042]);
module_output_bit_1043	m1043	(input_data_all[1796:0],output_data_all[1043]);
module_output_bit_1044	m1044	(input_data_all[1796:0],output_data_all[1044]);
module_output_bit_1045	m1045	(input_data_all[1796:0],output_data_all[1045]);
module_output_bit_1046	m1046	(input_data_all[1796:0],output_data_all[1046]);
module_output_bit_1047	m1047	(input_data_all[1796:0],output_data_all[1047]);
module_output_bit_1048	m1048	(input_data_all[1796:0],output_data_all[1048]);
module_output_bit_1049	m1049	(input_data_all[1796:0],output_data_all[1049]);
module_output_bit_1050	m1050	(input_data_all[1796:0],output_data_all[1050]);
module_output_bit_1051	m1051	(input_data_all[1796:0],output_data_all[1051]);
module_output_bit_1052	m1052	(input_data_all[1796:0],output_data_all[1052]);
module_output_bit_1053	m1053	(input_data_all[1796:0],output_data_all[1053]);
module_output_bit_1054	m1054	(input_data_all[1796:0],output_data_all[1054]);
module_output_bit_1055	m1055	(input_data_all[1796:0],output_data_all[1055]);
module_output_bit_1056	m1056	(input_data_all[1796:0],output_data_all[1056]);
module_output_bit_1057	m1057	(input_data_all[1796:0],output_data_all[1057]);
module_output_bit_1058	m1058	(input_data_all[1796:0],output_data_all[1058]);
module_output_bit_1059	m1059	(input_data_all[1796:0],output_data_all[1059]);
module_output_bit_1060	m1060	(input_data_all[1796:0],output_data_all[1060]);
module_output_bit_1061	m1061	(input_data_all[1796:0],output_data_all[1061]);
module_output_bit_1062	m1062	(input_data_all[1796:0],output_data_all[1062]);
module_output_bit_1063	m1063	(input_data_all[1796:0],output_data_all[1063]);
module_output_bit_1064	m1064	(input_data_all[1796:0],output_data_all[1064]);
module_output_bit_1065	m1065	(input_data_all[1796:0],output_data_all[1065]);
module_output_bit_1066	m1066	(input_data_all[1796:0],output_data_all[1066]);
module_output_bit_1067	m1067	(input_data_all[1796:0],output_data_all[1067]);
module_output_bit_1068	m1068	(input_data_all[1796:0],output_data_all[1068]);
module_output_bit_1069	m1069	(input_data_all[1796:0],output_data_all[1069]);
module_output_bit_1070	m1070	(input_data_all[1796:0],output_data_all[1070]);
module_output_bit_1071	m1071	(input_data_all[1796:0],output_data_all[1071]);
module_output_bit_1072	m1072	(input_data_all[1796:0],output_data_all[1072]);
module_output_bit_1073	m1073	(input_data_all[1796:0],output_data_all[1073]);
module_output_bit_1074	m1074	(input_data_all[1796:0],output_data_all[1074]);
module_output_bit_1075	m1075	(input_data_all[1796:0],output_data_all[1075]);
module_output_bit_1076	m1076	(input_data_all[1796:0],output_data_all[1076]);
module_output_bit_1077	m1077	(input_data_all[1796:0],output_data_all[1077]);
module_output_bit_1078	m1078	(input_data_all[1796:0],output_data_all[1078]);
module_output_bit_1079	m1079	(input_data_all[1796:0],output_data_all[1079]);
module_output_bit_1080	m1080	(input_data_all[1796:0],output_data_all[1080]);
module_output_bit_1081	m1081	(input_data_all[1796:0],output_data_all[1081]);
module_output_bit_1082	m1082	(input_data_all[1796:0],output_data_all[1082]);
module_output_bit_1083	m1083	(input_data_all[1796:0],output_data_all[1083]);
module_output_bit_1084	m1084	(input_data_all[1796:0],output_data_all[1084]);
module_output_bit_1085	m1085	(input_data_all[1796:0],output_data_all[1085]);
module_output_bit_1086	m1086	(input_data_all[1796:0],output_data_all[1086]);
module_output_bit_1087	m1087	(input_data_all[1796:0],output_data_all[1087]);
module_output_bit_1088	m1088	(input_data_all[1796:0],output_data_all[1088]);
module_output_bit_1089	m1089	(input_data_all[1796:0],output_data_all[1089]);
module_output_bit_1090	m1090	(input_data_all[1796:0],output_data_all[1090]);
module_output_bit_1091	m1091	(input_data_all[1796:0],output_data_all[1091]);
module_output_bit_1092	m1092	(input_data_all[1796:0],output_data_all[1092]);
module_output_bit_1093	m1093	(input_data_all[1796:0],output_data_all[1093]);
module_output_bit_1094	m1094	(input_data_all[1796:0],output_data_all[1094]);
module_output_bit_1095	m1095	(input_data_all[1796:0],output_data_all[1095]);
module_output_bit_1096	m1096	(input_data_all[1796:0],output_data_all[1096]);
module_output_bit_1097	m1097	(input_data_all[1796:0],output_data_all[1097]);
module_output_bit_1098	m1098	(input_data_all[1796:0],output_data_all[1098]);
module_output_bit_1099	m1099	(input_data_all[1796:0],output_data_all[1099]);
module_output_bit_1100	m1100	(input_data_all[1796:0],output_data_all[1100]);
module_output_bit_1101	m1101	(input_data_all[1796:0],output_data_all[1101]);
module_output_bit_1102	m1102	(input_data_all[1796:0],output_data_all[1102]);
module_output_bit_1103	m1103	(input_data_all[1796:0],output_data_all[1103]);
module_output_bit_1104	m1104	(input_data_all[1796:0],output_data_all[1104]);
module_output_bit_1105	m1105	(input_data_all[1796:0],output_data_all[1105]);
module_output_bit_1106	m1106	(input_data_all[1796:0],output_data_all[1106]);
module_output_bit_1107	m1107	(input_data_all[1796:0],output_data_all[1107]);
module_output_bit_1108	m1108	(input_data_all[1796:0],output_data_all[1108]);
module_output_bit_1109	m1109	(input_data_all[1796:0],output_data_all[1109]);
module_output_bit_1110	m1110	(input_data_all[1796:0],output_data_all[1110]);
module_output_bit_1111	m1111	(input_data_all[1796:0],output_data_all[1111]);
module_output_bit_1112	m1112	(input_data_all[1796:0],output_data_all[1112]);
module_output_bit_1113	m1113	(input_data_all[1796:0],output_data_all[1113]);
module_output_bit_1114	m1114	(input_data_all[1796:0],output_data_all[1114]);
module_output_bit_1115	m1115	(input_data_all[1796:0],output_data_all[1115]);
module_output_bit_1116	m1116	(input_data_all[1796:0],output_data_all[1116]);
module_output_bit_1117	m1117	(input_data_all[1796:0],output_data_all[1117]);
module_output_bit_1118	m1118	(input_data_all[1796:0],output_data_all[1118]);
module_output_bit_1119	m1119	(input_data_all[1796:0],output_data_all[1119]);
module_output_bit_1120	m1120	(input_data_all[1796:0],output_data_all[1120]);
module_output_bit_1121	m1121	(input_data_all[1796:0],output_data_all[1121]);
module_output_bit_1122	m1122	(input_data_all[1796:0],output_data_all[1122]);
module_output_bit_1123	m1123	(input_data_all[1796:0],output_data_all[1123]);
module_output_bit_1124	m1124	(input_data_all[1796:0],output_data_all[1124]);
module_output_bit_1125	m1125	(input_data_all[1796:0],output_data_all[1125]);
module_output_bit_1126	m1126	(input_data_all[1796:0],output_data_all[1126]);
module_output_bit_1127	m1127	(input_data_all[1796:0],output_data_all[1127]);
module_output_bit_1128	m1128	(input_data_all[1796:0],output_data_all[1128]);
module_output_bit_1129	m1129	(input_data_all[1796:0],output_data_all[1129]);
module_output_bit_1130	m1130	(input_data_all[1796:0],output_data_all[1130]);
module_output_bit_1131	m1131	(input_data_all[1796:0],output_data_all[1131]);
module_output_bit_1132	m1132	(input_data_all[1796:0],output_data_all[1132]);
module_output_bit_1133	m1133	(input_data_all[1796:0],output_data_all[1133]);
module_output_bit_1134	m1134	(input_data_all[1796:0],output_data_all[1134]);
module_output_bit_1135	m1135	(input_data_all[1796:0],output_data_all[1135]);
module_output_bit_1136	m1136	(input_data_all[1796:0],output_data_all[1136]);
module_output_bit_1137	m1137	(input_data_all[1796:0],output_data_all[1137]);
module_output_bit_1138	m1138	(input_data_all[1796:0],output_data_all[1138]);
module_output_bit_1139	m1139	(input_data_all[1796:0],output_data_all[1139]);
module_output_bit_1140	m1140	(input_data_all[1796:0],output_data_all[1140]);
module_output_bit_1141	m1141	(input_data_all[1796:0],output_data_all[1141]);
module_output_bit_1142	m1142	(input_data_all[1796:0],output_data_all[1142]);
module_output_bit_1143	m1143	(input_data_all[1796:0],output_data_all[1143]);
module_output_bit_1144	m1144	(input_data_all[1796:0],output_data_all[1144]);
module_output_bit_1145	m1145	(input_data_all[1796:0],output_data_all[1145]);
module_output_bit_1146	m1146	(input_data_all[1796:0],output_data_all[1146]);
module_output_bit_1147	m1147	(input_data_all[1796:0],output_data_all[1147]);
module_output_bit_1148	m1148	(input_data_all[1796:0],output_data_all[1148]);
module_output_bit_1149	m1149	(input_data_all[1796:0],output_data_all[1149]);
module_output_bit_1150	m1150	(input_data_all[1796:0],output_data_all[1150]);
module_output_bit_1151	m1151	(input_data_all[1796:0],output_data_all[1151]);
module_output_bit_1152	m1152	(input_data_all[1796:0],output_data_all[1152]);
module_output_bit_1153	m1153	(input_data_all[1796:0],output_data_all[1153]);
module_output_bit_1154	m1154	(input_data_all[1796:0],output_data_all[1154]);
module_output_bit_1155	m1155	(input_data_all[1796:0],output_data_all[1155]);
module_output_bit_1156	m1156	(input_data_all[1796:0],output_data_all[1156]);
module_output_bit_1157	m1157	(input_data_all[1796:0],output_data_all[1157]);
module_output_bit_1158	m1158	(input_data_all[1796:0],output_data_all[1158]);
module_output_bit_1159	m1159	(input_data_all[1796:0],output_data_all[1159]);
module_output_bit_1160	m1160	(input_data_all[1796:0],output_data_all[1160]);
module_output_bit_1161	m1161	(input_data_all[1796:0],output_data_all[1161]);
module_output_bit_1162	m1162	(input_data_all[1796:0],output_data_all[1162]);
module_output_bit_1163	m1163	(input_data_all[1796:0],output_data_all[1163]);
module_output_bit_1164	m1164	(input_data_all[1796:0],output_data_all[1164]);
module_output_bit_1165	m1165	(input_data_all[1796:0],output_data_all[1165]);
module_output_bit_1166	m1166	(input_data_all[1796:0],output_data_all[1166]);
module_output_bit_1167	m1167	(input_data_all[1796:0],output_data_all[1167]);
module_output_bit_1168	m1168	(input_data_all[1796:0],output_data_all[1168]);
module_output_bit_1169	m1169	(input_data_all[1796:0],output_data_all[1169]);
module_output_bit_1170	m1170	(input_data_all[1796:0],output_data_all[1170]);
module_output_bit_1171	m1171	(input_data_all[1796:0],output_data_all[1171]);
module_output_bit_1172	m1172	(input_data_all[1796:0],output_data_all[1172]);
module_output_bit_1173	m1173	(input_data_all[1796:0],output_data_all[1173]);
module_output_bit_1174	m1174	(input_data_all[1796:0],output_data_all[1174]);
module_output_bit_1175	m1175	(input_data_all[1796:0],output_data_all[1175]);
module_output_bit_1176	m1176	(input_data_all[1796:0],output_data_all[1176]);
module_output_bit_1177	m1177	(input_data_all[1796:0],output_data_all[1177]);
module_output_bit_1178	m1178	(input_data_all[1796:0],output_data_all[1178]);
module_output_bit_1179	m1179	(input_data_all[1796:0],output_data_all[1179]);
module_output_bit_1180	m1180	(input_data_all[1796:0],output_data_all[1180]);
module_output_bit_1181	m1181	(input_data_all[1796:0],output_data_all[1181]);
module_output_bit_1182	m1182	(input_data_all[1796:0],output_data_all[1182]);
module_output_bit_1183	m1183	(input_data_all[1796:0],output_data_all[1183]);
module_output_bit_1184	m1184	(input_data_all[1796:0],output_data_all[1184]);
module_output_bit_1185	m1185	(input_data_all[1796:0],output_data_all[1185]);
module_output_bit_1186	m1186	(input_data_all[1796:0],output_data_all[1186]);
module_output_bit_1187	m1187	(input_data_all[1796:0],output_data_all[1187]);
module_output_bit_1188	m1188	(input_data_all[1796:0],output_data_all[1188]);
module_output_bit_1189	m1189	(input_data_all[1796:0],output_data_all[1189]);
module_output_bit_1190	m1190	(input_data_all[1796:0],output_data_all[1190]);
module_output_bit_1191	m1191	(input_data_all[1796:0],output_data_all[1191]);
module_output_bit_1192	m1192	(input_data_all[1796:0],output_data_all[1192]);
module_output_bit_1193	m1193	(input_data_all[1796:0],output_data_all[1193]);
module_output_bit_1194	m1194	(input_data_all[1796:0],output_data_all[1194]);
module_output_bit_1195	m1195	(input_data_all[1796:0],output_data_all[1195]);
module_output_bit_1196	m1196	(input_data_all[1796:0],output_data_all[1196]);
module_output_bit_1197	m1197	(input_data_all[1796:0],output_data_all[1197]);
module_output_bit_1198	m1198	(input_data_all[1796:0],output_data_all[1198]);
module_output_bit_1199	m1199	(input_data_all[1796:0],output_data_all[1199]);
module_output_bit_1200	m1200	(input_data_all[1796:0],output_data_all[1200]);
module_output_bit_1201	m1201	(input_data_all[1796:0],output_data_all[1201]);
module_output_bit_1202	m1202	(input_data_all[1796:0],output_data_all[1202]);
module_output_bit_1203	m1203	(input_data_all[1796:0],output_data_all[1203]);
module_output_bit_1204	m1204	(input_data_all[1796:0],output_data_all[1204]);
module_output_bit_1205	m1205	(input_data_all[1796:0],output_data_all[1205]);
module_output_bit_1206	m1206	(input_data_all[1796:0],output_data_all[1206]);
module_output_bit_1207	m1207	(input_data_all[1796:0],output_data_all[1207]);
module_output_bit_1208	m1208	(input_data_all[1796:0],output_data_all[1208]);
module_output_bit_1209	m1209	(input_data_all[1796:0],output_data_all[1209]);
module_output_bit_1210	m1210	(input_data_all[1796:0],output_data_all[1210]);
module_output_bit_1211	m1211	(input_data_all[1796:0],output_data_all[1211]);
module_output_bit_1212	m1212	(input_data_all[1796:0],output_data_all[1212]);
module_output_bit_1213	m1213	(input_data_all[1796:0],output_data_all[1213]);
module_output_bit_1214	m1214	(input_data_all[1796:0],output_data_all[1214]);
module_output_bit_1215	m1215	(input_data_all[1796:0],output_data_all[1215]);
module_output_bit_1216	m1216	(input_data_all[1796:0],output_data_all[1216]);
module_output_bit_1217	m1217	(input_data_all[1796:0],output_data_all[1217]);
module_output_bit_1218	m1218	(input_data_all[1796:0],output_data_all[1218]);
module_output_bit_1219	m1219	(input_data_all[1796:0],output_data_all[1219]);
module_output_bit_1220	m1220	(input_data_all[1796:0],output_data_all[1220]);
module_output_bit_1221	m1221	(input_data_all[1796:0],output_data_all[1221]);
module_output_bit_1222	m1222	(input_data_all[1796:0],output_data_all[1222]);
module_output_bit_1223	m1223	(input_data_all[1796:0],output_data_all[1223]);
module_output_bit_1224	m1224	(input_data_all[1796:0],output_data_all[1224]);
module_output_bit_1225	m1225	(input_data_all[1796:0],output_data_all[1225]);
module_output_bit_1226	m1226	(input_data_all[1796:0],output_data_all[1226]);
module_output_bit_1227	m1227	(input_data_all[1796:0],output_data_all[1227]);
module_output_bit_1228	m1228	(input_data_all[1796:0],output_data_all[1228]);
module_output_bit_1229	m1229	(input_data_all[1796:0],output_data_all[1229]);
module_output_bit_1230	m1230	(input_data_all[1796:0],output_data_all[1230]);
module_output_bit_1231	m1231	(input_data_all[1796:0],output_data_all[1231]);
module_output_bit_1232	m1232	(input_data_all[1796:0],output_data_all[1232]);
module_output_bit_1233	m1233	(input_data_all[1796:0],output_data_all[1233]);
module_output_bit_1234	m1234	(input_data_all[1796:0],output_data_all[1234]);
module_output_bit_1235	m1235	(input_data_all[1796:0],output_data_all[1235]);
module_output_bit_1236	m1236	(input_data_all[1796:0],output_data_all[1236]);
module_output_bit_1237	m1237	(input_data_all[1796:0],output_data_all[1237]);
module_output_bit_1238	m1238	(input_data_all[1796:0],output_data_all[1238]);
module_output_bit_1239	m1239	(input_data_all[1796:0],output_data_all[1239]);
module_output_bit_1240	m1240	(input_data_all[1796:0],output_data_all[1240]);
module_output_bit_1241	m1241	(input_data_all[1796:0],output_data_all[1241]);
module_output_bit_1242	m1242	(input_data_all[1796:0],output_data_all[1242]);
module_output_bit_1243	m1243	(input_data_all[1796:0],output_data_all[1243]);
module_output_bit_1244	m1244	(input_data_all[1796:0],output_data_all[1244]);
module_output_bit_1245	m1245	(input_data_all[1796:0],output_data_all[1245]);
module_output_bit_1246	m1246	(input_data_all[1796:0],output_data_all[1246]);
module_output_bit_1247	m1247	(input_data_all[1796:0],output_data_all[1247]);
module_output_bit_1248	m1248	(input_data_all[1796:0],output_data_all[1248]);
module_output_bit_1249	m1249	(input_data_all[1796:0],output_data_all[1249]);
module_output_bit_1250	m1250	(input_data_all[1796:0],output_data_all[1250]);
module_output_bit_1251	m1251	(input_data_all[1796:0],output_data_all[1251]);
module_output_bit_1252	m1252	(input_data_all[1796:0],output_data_all[1252]);
module_output_bit_1253	m1253	(input_data_all[1796:0],output_data_all[1253]);
module_output_bit_1254	m1254	(input_data_all[1796:0],output_data_all[1254]);
module_output_bit_1255	m1255	(input_data_all[1796:0],output_data_all[1255]);
module_output_bit_1256	m1256	(input_data_all[1796:0],output_data_all[1256]);
module_output_bit_1257	m1257	(input_data_all[1796:0],output_data_all[1257]);
module_output_bit_1258	m1258	(input_data_all[1796:0],output_data_all[1258]);
module_output_bit_1259	m1259	(input_data_all[1796:0],output_data_all[1259]);
module_output_bit_1260	m1260	(input_data_all[1796:0],output_data_all[1260]);
module_output_bit_1261	m1261	(input_data_all[1796:0],output_data_all[1261]);
module_output_bit_1262	m1262	(input_data_all[1796:0],output_data_all[1262]);
module_output_bit_1263	m1263	(input_data_all[1796:0],output_data_all[1263]);
module_output_bit_1264	m1264	(input_data_all[1796:0],output_data_all[1264]);
module_output_bit_1265	m1265	(input_data_all[1796:0],output_data_all[1265]);
module_output_bit_1266	m1266	(input_data_all[1796:0],output_data_all[1266]);
module_output_bit_1267	m1267	(input_data_all[1796:0],output_data_all[1267]);
module_output_bit_1268	m1268	(input_data_all[1796:0],output_data_all[1268]);
module_output_bit_1269	m1269	(input_data_all[1796:0],output_data_all[1269]);
module_output_bit_1270	m1270	(input_data_all[1796:0],output_data_all[1270]);
module_output_bit_1271	m1271	(input_data_all[1796:0],output_data_all[1271]);
module_output_bit_1272	m1272	(input_data_all[1796:0],output_data_all[1272]);
module_output_bit_1273	m1273	(input_data_all[1796:0],output_data_all[1273]);
module_output_bit_1274	m1274	(input_data_all[1796:0],output_data_all[1274]);
module_output_bit_1275	m1275	(input_data_all[1796:0],output_data_all[1275]);
module_output_bit_1276	m1276	(input_data_all[1796:0],output_data_all[1276]);
module_output_bit_1277	m1277	(input_data_all[1796:0],output_data_all[1277]);
module_output_bit_1278	m1278	(input_data_all[1796:0],output_data_all[1278]);
module_output_bit_1279	m1279	(input_data_all[1796:0],output_data_all[1279]);
module_output_bit_1280	m1280	(input_data_all[1796:0],output_data_all[1280]);
module_output_bit_1281	m1281	(input_data_all[1796:0],output_data_all[1281]);
module_output_bit_1282	m1282	(input_data_all[1796:0],output_data_all[1282]);
module_output_bit_1283	m1283	(input_data_all[1796:0],output_data_all[1283]);
module_output_bit_1284	m1284	(input_data_all[1796:0],output_data_all[1284]);
module_output_bit_1285	m1285	(input_data_all[1796:0],output_data_all[1285]);
module_output_bit_1286	m1286	(input_data_all[1796:0],output_data_all[1286]);
module_output_bit_1287	m1287	(input_data_all[1796:0],output_data_all[1287]);
module_output_bit_1288	m1288	(input_data_all[1796:0],output_data_all[1288]);
module_output_bit_1289	m1289	(input_data_all[1796:0],output_data_all[1289]);
module_output_bit_1290	m1290	(input_data_all[1796:0],output_data_all[1290]);
module_output_bit_1291	m1291	(input_data_all[1796:0],output_data_all[1291]);
module_output_bit_1292	m1292	(input_data_all[1796:0],output_data_all[1292]);
module_output_bit_1293	m1293	(input_data_all[1796:0],output_data_all[1293]);
module_output_bit_1294	m1294	(input_data_all[1796:0],output_data_all[1294]);
module_output_bit_1295	m1295	(input_data_all[1796:0],output_data_all[1295]);
module_output_bit_1296	m1296	(input_data_all[1796:0],output_data_all[1296]);
module_output_bit_1297	m1297	(input_data_all[1796:0],output_data_all[1297]);
module_output_bit_1298	m1298	(input_data_all[1796:0],output_data_all[1298]);
module_output_bit_1299	m1299	(input_data_all[1796:0],output_data_all[1299]);
module_output_bit_1300	m1300	(input_data_all[1796:0],output_data_all[1300]);
module_output_bit_1301	m1301	(input_data_all[1796:0],output_data_all[1301]);
module_output_bit_1302	m1302	(input_data_all[1796:0],output_data_all[1302]);
module_output_bit_1303	m1303	(input_data_all[1796:0],output_data_all[1303]);
module_output_bit_1304	m1304	(input_data_all[1796:0],output_data_all[1304]);
module_output_bit_1305	m1305	(input_data_all[1796:0],output_data_all[1305]);
module_output_bit_1306	m1306	(input_data_all[1796:0],output_data_all[1306]);
module_output_bit_1307	m1307	(input_data_all[1796:0],output_data_all[1307]);
module_output_bit_1308	m1308	(input_data_all[1796:0],output_data_all[1308]);
module_output_bit_1309	m1309	(input_data_all[1796:0],output_data_all[1309]);
module_output_bit_1310	m1310	(input_data_all[1796:0],output_data_all[1310]);
module_output_bit_1311	m1311	(input_data_all[1796:0],output_data_all[1311]);
module_output_bit_1312	m1312	(input_data_all[1796:0],output_data_all[1312]);
module_output_bit_1313	m1313	(input_data_all[1796:0],output_data_all[1313]);
module_output_bit_1314	m1314	(input_data_all[1796:0],output_data_all[1314]);
module_output_bit_1315	m1315	(input_data_all[1796:0],output_data_all[1315]);
module_output_bit_1316	m1316	(input_data_all[1796:0],output_data_all[1316]);
module_output_bit_1317	m1317	(input_data_all[1796:0],output_data_all[1317]);
module_output_bit_1318	m1318	(input_data_all[1796:0],output_data_all[1318]);
module_output_bit_1319	m1319	(input_data_all[1796:0],output_data_all[1319]);
module_output_bit_1320	m1320	(input_data_all[1796:0],output_data_all[1320]);
module_output_bit_1321	m1321	(input_data_all[1796:0],output_data_all[1321]);
module_output_bit_1322	m1322	(input_data_all[1796:0],output_data_all[1322]);
module_output_bit_1323	m1323	(input_data_all[1796:0],output_data_all[1323]);
module_output_bit_1324	m1324	(input_data_all[1796:0],output_data_all[1324]);
module_output_bit_1325	m1325	(input_data_all[1796:0],output_data_all[1325]);
module_output_bit_1326	m1326	(input_data_all[1796:0],output_data_all[1326]);
module_output_bit_1327	m1327	(input_data_all[1796:0],output_data_all[1327]);
module_output_bit_1328	m1328	(input_data_all[1796:0],output_data_all[1328]);
module_output_bit_1329	m1329	(input_data_all[1796:0],output_data_all[1329]);
module_output_bit_1330	m1330	(input_data_all[1796:0],output_data_all[1330]);
module_output_bit_1331	m1331	(input_data_all[1796:0],output_data_all[1331]);
module_output_bit_1332	m1332	(input_data_all[1796:0],output_data_all[1332]);
module_output_bit_1333	m1333	(input_data_all[1796:0],output_data_all[1333]);
module_output_bit_1334	m1334	(input_data_all[1796:0],output_data_all[1334]);
module_output_bit_1335	m1335	(input_data_all[1796:0],output_data_all[1335]);
module_output_bit_1336	m1336	(input_data_all[1796:0],output_data_all[1336]);
module_output_bit_1337	m1337	(input_data_all[1796:0],output_data_all[1337]);
module_output_bit_1338	m1338	(input_data_all[1796:0],output_data_all[1338]);
module_output_bit_1339	m1339	(input_data_all[1796:0],output_data_all[1339]);
module_output_bit_1340	m1340	(input_data_all[1796:0],output_data_all[1340]);
module_output_bit_1341	m1341	(input_data_all[1796:0],output_data_all[1341]);
module_output_bit_1342	m1342	(input_data_all[1796:0],output_data_all[1342]);
module_output_bit_1343	m1343	(input_data_all[1796:0],output_data_all[1343]);
module_output_bit_1344	m1344	(input_data_all[1796:0],output_data_all[1344]);
module_output_bit_1345	m1345	(input_data_all[1796:0],output_data_all[1345]);
module_output_bit_1346	m1346	(input_data_all[1796:0],output_data_all[1346]);
module_output_bit_1347	m1347	(input_data_all[1796:0],output_data_all[1347]);
module_output_bit_1348	m1348	(input_data_all[1796:0],output_data_all[1348]);
module_output_bit_1349	m1349	(input_data_all[1796:0],output_data_all[1349]);
module_output_bit_1350	m1350	(input_data_all[1796:0],output_data_all[1350]);
module_output_bit_1351	m1351	(input_data_all[1796:0],output_data_all[1351]);
module_output_bit_1352	m1352	(input_data_all[1796:0],output_data_all[1352]);
module_output_bit_1353	m1353	(input_data_all[1796:0],output_data_all[1353]);
module_output_bit_1354	m1354	(input_data_all[1796:0],output_data_all[1354]);
module_output_bit_1355	m1355	(input_data_all[1796:0],output_data_all[1355]);
module_output_bit_1356	m1356	(input_data_all[1796:0],output_data_all[1356]);
module_output_bit_1357	m1357	(input_data_all[1796:0],output_data_all[1357]);
module_output_bit_1358	m1358	(input_data_all[1796:0],output_data_all[1358]);
module_output_bit_1359	m1359	(input_data_all[1796:0],output_data_all[1359]);
module_output_bit_1360	m1360	(input_data_all[1796:0],output_data_all[1360]);
module_output_bit_1361	m1361	(input_data_all[1796:0],output_data_all[1361]);
module_output_bit_1362	m1362	(input_data_all[1796:0],output_data_all[1362]);
module_output_bit_1363	m1363	(input_data_all[1796:0],output_data_all[1363]);
module_output_bit_1364	m1364	(input_data_all[1796:0],output_data_all[1364]);
module_output_bit_1365	m1365	(input_data_all[1796:0],output_data_all[1365]);
module_output_bit_1366	m1366	(input_data_all[1796:0],output_data_all[1366]);
module_output_bit_1367	m1367	(input_data_all[1796:0],output_data_all[1367]);
module_output_bit_1368	m1368	(input_data_all[1796:0],output_data_all[1368]);
module_output_bit_1369	m1369	(input_data_all[1796:0],output_data_all[1369]);
module_output_bit_1370	m1370	(input_data_all[1796:0],output_data_all[1370]);
module_output_bit_1371	m1371	(input_data_all[1796:0],output_data_all[1371]);
module_output_bit_1372	m1372	(input_data_all[1796:0],output_data_all[1372]);
module_output_bit_1373	m1373	(input_data_all[1796:0],output_data_all[1373]);
module_output_bit_1374	m1374	(input_data_all[1796:0],output_data_all[1374]);
module_output_bit_1375	m1375	(input_data_all[1796:0],output_data_all[1375]);
module_output_bit_1376	m1376	(input_data_all[1796:0],output_data_all[1376]);
module_output_bit_1377	m1377	(input_data_all[1796:0],output_data_all[1377]);
module_output_bit_1378	m1378	(input_data_all[1796:0],output_data_all[1378]);
module_output_bit_1379	m1379	(input_data_all[1796:0],output_data_all[1379]);
module_output_bit_1380	m1380	(input_data_all[1796:0],output_data_all[1380]);
module_output_bit_1381	m1381	(input_data_all[1796:0],output_data_all[1381]);
module_output_bit_1382	m1382	(input_data_all[1796:0],output_data_all[1382]);
module_output_bit_1383	m1383	(input_data_all[1796:0],output_data_all[1383]);
module_output_bit_1384	m1384	(input_data_all[1796:0],output_data_all[1384]);
module_output_bit_1385	m1385	(input_data_all[1796:0],output_data_all[1385]);
module_output_bit_1386	m1386	(input_data_all[1796:0],output_data_all[1386]);
module_output_bit_1387	m1387	(input_data_all[1796:0],output_data_all[1387]);
module_output_bit_1388	m1388	(input_data_all[1796:0],output_data_all[1388]);
module_output_bit_1389	m1389	(input_data_all[1796:0],output_data_all[1389]);
module_output_bit_1390	m1390	(input_data_all[1796:0],output_data_all[1390]);
module_output_bit_1391	m1391	(input_data_all[1796:0],output_data_all[1391]);
module_output_bit_1392	m1392	(input_data_all[1796:0],output_data_all[1392]);
module_output_bit_1393	m1393	(input_data_all[1796:0],output_data_all[1393]);
module_output_bit_1394	m1394	(input_data_all[1796:0],output_data_all[1394]);
module_output_bit_1395	m1395	(input_data_all[1796:0],output_data_all[1395]);
module_output_bit_1396	m1396	(input_data_all[1796:0],output_data_all[1396]);
module_output_bit_1397	m1397	(input_data_all[1796:0],output_data_all[1397]);
module_output_bit_1398	m1398	(input_data_all[1796:0],output_data_all[1398]);
module_output_bit_1399	m1399	(input_data_all[1796:0],output_data_all[1399]);
module_output_bit_1400	m1400	(input_data_all[1796:0],output_data_all[1400]);
module_output_bit_1401	m1401	(input_data_all[1796:0],output_data_all[1401]);
module_output_bit_1402	m1402	(input_data_all[1796:0],output_data_all[1402]);
module_output_bit_1403	m1403	(input_data_all[1796:0],output_data_all[1403]);
module_output_bit_1404	m1404	(input_data_all[1796:0],output_data_all[1404]);
module_output_bit_1405	m1405	(input_data_all[1796:0],output_data_all[1405]);
module_output_bit_1406	m1406	(input_data_all[1796:0],output_data_all[1406]);
module_output_bit_1407	m1407	(input_data_all[1796:0],output_data_all[1407]);
module_output_bit_1408	m1408	(input_data_all[1796:0],output_data_all[1408]);
module_output_bit_1409	m1409	(input_data_all[1796:0],output_data_all[1409]);
module_output_bit_1410	m1410	(input_data_all[1796:0],output_data_all[1410]);
module_output_bit_1411	m1411	(input_data_all[1796:0],output_data_all[1411]);
module_output_bit_1412	m1412	(input_data_all[1796:0],output_data_all[1412]);
module_output_bit_1413	m1413	(input_data_all[1796:0],output_data_all[1413]);
module_output_bit_1414	m1414	(input_data_all[1796:0],output_data_all[1414]);
module_output_bit_1415	m1415	(input_data_all[1796:0],output_data_all[1415]);
module_output_bit_1416	m1416	(input_data_all[1796:0],output_data_all[1416]);
module_output_bit_1417	m1417	(input_data_all[1796:0],output_data_all[1417]);
module_output_bit_1418	m1418	(input_data_all[1796:0],output_data_all[1418]);
module_output_bit_1419	m1419	(input_data_all[1796:0],output_data_all[1419]);
module_output_bit_1420	m1420	(input_data_all[1796:0],output_data_all[1420]);
module_output_bit_1421	m1421	(input_data_all[1796:0],output_data_all[1421]);
module_output_bit_1422	m1422	(input_data_all[1796:0],output_data_all[1422]);
module_output_bit_1423	m1423	(input_data_all[1796:0],output_data_all[1423]);
module_output_bit_1424	m1424	(input_data_all[1796:0],output_data_all[1424]);
module_output_bit_1425	m1425	(input_data_all[1796:0],output_data_all[1425]);
module_output_bit_1426	m1426	(input_data_all[1796:0],output_data_all[1426]);
module_output_bit_1427	m1427	(input_data_all[1796:0],output_data_all[1427]);
module_output_bit_1428	m1428	(input_data_all[1796:0],output_data_all[1428]);
module_output_bit_1429	m1429	(input_data_all[1796:0],output_data_all[1429]);
module_output_bit_1430	m1430	(input_data_all[1796:0],output_data_all[1430]);
module_output_bit_1431	m1431	(input_data_all[1796:0],output_data_all[1431]);
module_output_bit_1432	m1432	(input_data_all[1796:0],output_data_all[1432]);
module_output_bit_1433	m1433	(input_data_all[1796:0],output_data_all[1433]);
module_output_bit_1434	m1434	(input_data_all[1796:0],output_data_all[1434]);
module_output_bit_1435	m1435	(input_data_all[1796:0],output_data_all[1435]);
module_output_bit_1436	m1436	(input_data_all[1796:0],output_data_all[1436]);
module_output_bit_1437	m1437	(input_data_all[1796:0],output_data_all[1437]);
module_output_bit_1438	m1438	(input_data_all[1796:0],output_data_all[1438]);
module_output_bit_1439	m1439	(input_data_all[1796:0],output_data_all[1439]);
module_output_bit_1440	m1440	(input_data_all[1796:0],output_data_all[1440]);
module_output_bit_1441	m1441	(input_data_all[1796:0],output_data_all[1441]);
module_output_bit_1442	m1442	(input_data_all[1796:0],output_data_all[1442]);
module_output_bit_1443	m1443	(input_data_all[1796:0],output_data_all[1443]);
module_output_bit_1444	m1444	(input_data_all[1796:0],output_data_all[1444]);
module_output_bit_1445	m1445	(input_data_all[1796:0],output_data_all[1445]);
module_output_bit_1446	m1446	(input_data_all[1796:0],output_data_all[1446]);
module_output_bit_1447	m1447	(input_data_all[1796:0],output_data_all[1447]);
module_output_bit_1448	m1448	(input_data_all[1796:0],output_data_all[1448]);
module_output_bit_1449	m1449	(input_data_all[1796:0],output_data_all[1449]);
module_output_bit_1450	m1450	(input_data_all[1796:0],output_data_all[1450]);
module_output_bit_1451	m1451	(input_data_all[1796:0],output_data_all[1451]);
module_output_bit_1452	m1452	(input_data_all[1796:0],output_data_all[1452]);
module_output_bit_1453	m1453	(input_data_all[1796:0],output_data_all[1453]);
module_output_bit_1454	m1454	(input_data_all[1796:0],output_data_all[1454]);
module_output_bit_1455	m1455	(input_data_all[1796:0],output_data_all[1455]);
module_output_bit_1456	m1456	(input_data_all[1796:0],output_data_all[1456]);
module_output_bit_1457	m1457	(input_data_all[1796:0],output_data_all[1457]);
module_output_bit_1458	m1458	(input_data_all[1796:0],output_data_all[1458]);
module_output_bit_1459	m1459	(input_data_all[1796:0],output_data_all[1459]);
module_output_bit_1460	m1460	(input_data_all[1796:0],output_data_all[1460]);
module_output_bit_1461	m1461	(input_data_all[1796:0],output_data_all[1461]);
module_output_bit_1462	m1462	(input_data_all[1796:0],output_data_all[1462]);
module_output_bit_1463	m1463	(input_data_all[1796:0],output_data_all[1463]);
module_output_bit_1464	m1464	(input_data_all[1796:0],output_data_all[1464]);
module_output_bit_1465	m1465	(input_data_all[1796:0],output_data_all[1465]);
module_output_bit_1466	m1466	(input_data_all[1796:0],output_data_all[1466]);
module_output_bit_1467	m1467	(input_data_all[1796:0],output_data_all[1467]);
module_output_bit_1468	m1468	(input_data_all[1796:0],output_data_all[1468]);
module_output_bit_1469	m1469	(input_data_all[1796:0],output_data_all[1469]);
module_output_bit_1470	m1470	(input_data_all[1796:0],output_data_all[1470]);
module_output_bit_1471	m1471	(input_data_all[1796:0],output_data_all[1471]);
module_output_bit_1472	m1472	(input_data_all[1796:0],output_data_all[1472]);
module_output_bit_1473	m1473	(input_data_all[1796:0],output_data_all[1473]);
module_output_bit_1474	m1474	(input_data_all[1796:0],output_data_all[1474]);
module_output_bit_1475	m1475	(input_data_all[1796:0],output_data_all[1475]);
module_output_bit_1476	m1476	(input_data_all[1796:0],output_data_all[1476]);
module_output_bit_1477	m1477	(input_data_all[1796:0],output_data_all[1477]);
module_output_bit_1478	m1478	(input_data_all[1796:0],output_data_all[1478]);
module_output_bit_1479	m1479	(input_data_all[1796:0],output_data_all[1479]);
module_output_bit_1480	m1480	(input_data_all[1796:0],output_data_all[1480]);
module_output_bit_1481	m1481	(input_data_all[1796:0],output_data_all[1481]);
module_output_bit_1482	m1482	(input_data_all[1796:0],output_data_all[1482]);
module_output_bit_1483	m1483	(input_data_all[1796:0],output_data_all[1483]);
module_output_bit_1484	m1484	(input_data_all[1796:0],output_data_all[1484]);
module_output_bit_1485	m1485	(input_data_all[1796:0],output_data_all[1485]);
module_output_bit_1486	m1486	(input_data_all[1796:0],output_data_all[1486]);
module_output_bit_1487	m1487	(input_data_all[1796:0],output_data_all[1487]);
module_output_bit_1488	m1488	(input_data_all[1796:0],output_data_all[1488]);
module_output_bit_1489	m1489	(input_data_all[1796:0],output_data_all[1489]);
module_output_bit_1490	m1490	(input_data_all[1796:0],output_data_all[1490]);
module_output_bit_1491	m1491	(input_data_all[1796:0],output_data_all[1491]);
module_output_bit_1492	m1492	(input_data_all[1796:0],output_data_all[1492]);
module_output_bit_1493	m1493	(input_data_all[1796:0],output_data_all[1493]);
module_output_bit_1494	m1494	(input_data_all[1796:0],output_data_all[1494]);
module_output_bit_1495	m1495	(input_data_all[1796:0],output_data_all[1495]);
module_output_bit_1496	m1496	(input_data_all[1796:0],output_data_all[1496]);
module_output_bit_1497	m1497	(input_data_all[1796:0],output_data_all[1497]);
module_output_bit_1498	m1498	(input_data_all[1796:0],output_data_all[1498]);
module_output_bit_1499	m1499	(input_data_all[1796:0],output_data_all[1499]);
module_output_bit_1500	m1500	(input_data_all[1796:0],output_data_all[1500]);
module_output_bit_1501	m1501	(input_data_all[1796:0],output_data_all[1501]);
module_output_bit_1502	m1502	(input_data_all[1796:0],output_data_all[1502]);
module_output_bit_1503	m1503	(input_data_all[1796:0],output_data_all[1503]);
module_output_bit_1504	m1504	(input_data_all[1796:0],output_data_all[1504]);
module_output_bit_1505	m1505	(input_data_all[1796:0],output_data_all[1505]);
module_output_bit_1506	m1506	(input_data_all[1796:0],output_data_all[1506]);
module_output_bit_1507	m1507	(input_data_all[1796:0],output_data_all[1507]);
module_output_bit_1508	m1508	(input_data_all[1796:0],output_data_all[1508]);
module_output_bit_1509	m1509	(input_data_all[1796:0],output_data_all[1509]);
module_output_bit_1510	m1510	(input_data_all[1796:0],output_data_all[1510]);
module_output_bit_1511	m1511	(input_data_all[1796:0],output_data_all[1511]);
module_output_bit_1512	m1512	(input_data_all[1796:0],output_data_all[1512]);
module_output_bit_1513	m1513	(input_data_all[1796:0],output_data_all[1513]);
module_output_bit_1514	m1514	(input_data_all[1796:0],output_data_all[1514]);
module_output_bit_1515	m1515	(input_data_all[1796:0],output_data_all[1515]);
module_output_bit_1516	m1516	(input_data_all[1796:0],output_data_all[1516]);
module_output_bit_1517	m1517	(input_data_all[1796:0],output_data_all[1517]);
module_output_bit_1518	m1518	(input_data_all[1796:0],output_data_all[1518]);
module_output_bit_1519	m1519	(input_data_all[1796:0],output_data_all[1519]);
module_output_bit_1520	m1520	(input_data_all[1796:0],output_data_all[1520]);
module_output_bit_1521	m1521	(input_data_all[1796:0],output_data_all[1521]);
module_output_bit_1522	m1522	(input_data_all[1796:0],output_data_all[1522]);
module_output_bit_1523	m1523	(input_data_all[1796:0],output_data_all[1523]);
module_output_bit_1524	m1524	(input_data_all[1796:0],output_data_all[1524]);
module_output_bit_1525	m1525	(input_data_all[1796:0],output_data_all[1525]);
module_output_bit_1526	m1526	(input_data_all[1796:0],output_data_all[1526]);
module_output_bit_1527	m1527	(input_data_all[1796:0],output_data_all[1527]);
module_output_bit_1528	m1528	(input_data_all[1796:0],output_data_all[1528]);
module_output_bit_1529	m1529	(input_data_all[1796:0],output_data_all[1529]);
module_output_bit_1530	m1530	(input_data_all[1796:0],output_data_all[1530]);
module_output_bit_1531	m1531	(input_data_all[1796:0],output_data_all[1531]);
module_output_bit_1532	m1532	(input_data_all[1796:0],output_data_all[1532]);
module_output_bit_1533	m1533	(input_data_all[1796:0],output_data_all[1533]);
module_output_bit_1534	m1534	(input_data_all[1796:0],output_data_all[1534]);
module_output_bit_1535	m1535	(input_data_all[1796:0],output_data_all[1535]);
module_output_bit_1536	m1536	(input_data_all[1796:0],output_data_all[1536]);
module_output_bit_1537	m1537	(input_data_all[1796:0],output_data_all[1537]);
module_output_bit_1538	m1538	(input_data_all[1796:0],output_data_all[1538]);
module_output_bit_1539	m1539	(input_data_all[1796:0],output_data_all[1539]);
module_output_bit_1540	m1540	(input_data_all[1796:0],output_data_all[1540]);
module_output_bit_1541	m1541	(input_data_all[1796:0],output_data_all[1541]);
module_output_bit_1542	m1542	(input_data_all[1796:0],output_data_all[1542]);
module_output_bit_1543	m1543	(input_data_all[1796:0],output_data_all[1543]);
module_output_bit_1544	m1544	(input_data_all[1796:0],output_data_all[1544]);
module_output_bit_1545	m1545	(input_data_all[1796:0],output_data_all[1545]);
module_output_bit_1546	m1546	(input_data_all[1796:0],output_data_all[1546]);
module_output_bit_1547	m1547	(input_data_all[1796:0],output_data_all[1547]);
module_output_bit_1548	m1548	(input_data_all[1796:0],output_data_all[1548]);
module_output_bit_1549	m1549	(input_data_all[1796:0],output_data_all[1549]);
module_output_bit_1550	m1550	(input_data_all[1796:0],output_data_all[1550]);
module_output_bit_1551	m1551	(input_data_all[1796:0],output_data_all[1551]);
module_output_bit_1552	m1552	(input_data_all[1796:0],output_data_all[1552]);
module_output_bit_1553	m1553	(input_data_all[1796:0],output_data_all[1553]);
module_output_bit_1554	m1554	(input_data_all[1796:0],output_data_all[1554]);
module_output_bit_1555	m1555	(input_data_all[1796:0],output_data_all[1555]);
module_output_bit_1556	m1556	(input_data_all[1796:0],output_data_all[1556]);
module_output_bit_1557	m1557	(input_data_all[1796:0],output_data_all[1557]);
module_output_bit_1558	m1558	(input_data_all[1796:0],output_data_all[1558]);
module_output_bit_1559	m1559	(input_data_all[1796:0],output_data_all[1559]);
module_output_bit_1560	m1560	(input_data_all[1796:0],output_data_all[1560]);
module_output_bit_1561	m1561	(input_data_all[1796:0],output_data_all[1561]);
module_output_bit_1562	m1562	(input_data_all[1796:0],output_data_all[1562]);
module_output_bit_1563	m1563	(input_data_all[1796:0],output_data_all[1563]);
module_output_bit_1564	m1564	(input_data_all[1796:0],output_data_all[1564]);
module_output_bit_1565	m1565	(input_data_all[1796:0],output_data_all[1565]);
module_output_bit_1566	m1566	(input_data_all[1796:0],output_data_all[1566]);
module_output_bit_1567	m1567	(input_data_all[1796:0],output_data_all[1567]);
module_output_bit_1568	m1568	(input_data_all[1796:0],output_data_all[1568]);
module_output_bit_1569	m1569	(input_data_all[1796:0],output_data_all[1569]);
module_output_bit_1570	m1570	(input_data_all[1796:0],output_data_all[1570]);
module_output_bit_1571	m1571	(input_data_all[1796:0],output_data_all[1571]);
module_output_bit_1572	m1572	(input_data_all[1796:0],output_data_all[1572]);
module_output_bit_1573	m1573	(input_data_all[1796:0],output_data_all[1573]);
module_output_bit_1574	m1574	(input_data_all[1796:0],output_data_all[1574]);
module_output_bit_1575	m1575	(input_data_all[1796:0],output_data_all[1575]);
module_output_bit_1576	m1576	(input_data_all[1796:0],output_data_all[1576]);
module_output_bit_1577	m1577	(input_data_all[1796:0],output_data_all[1577]);
module_output_bit_1578	m1578	(input_data_all[1796:0],output_data_all[1578]);
module_output_bit_1579	m1579	(input_data_all[1796:0],output_data_all[1579]);
module_output_bit_1580	m1580	(input_data_all[1796:0],output_data_all[1580]);
module_output_bit_1581	m1581	(input_data_all[1796:0],output_data_all[1581]);
module_output_bit_1582	m1582	(input_data_all[1796:0],output_data_all[1582]);
module_output_bit_1583	m1583	(input_data_all[1796:0],output_data_all[1583]);
module_output_bit_1584	m1584	(input_data_all[1796:0],output_data_all[1584]);
module_output_bit_1585	m1585	(input_data_all[1796:0],output_data_all[1585]);
module_output_bit_1586	m1586	(input_data_all[1796:0],output_data_all[1586]);
module_output_bit_1587	m1587	(input_data_all[1796:0],output_data_all[1587]);
module_output_bit_1588	m1588	(input_data_all[1796:0],output_data_all[1588]);
module_output_bit_1589	m1589	(input_data_all[1796:0],output_data_all[1589]);
module_output_bit_1590	m1590	(input_data_all[1796:0],output_data_all[1590]);
module_output_bit_1591	m1591	(input_data_all[1796:0],output_data_all[1591]);
module_output_bit_1592	m1592	(input_data_all[1796:0],output_data_all[1592]);
module_output_bit_1593	m1593	(input_data_all[1796:0],output_data_all[1593]);
module_output_bit_1594	m1594	(input_data_all[1796:0],output_data_all[1594]);
module_output_bit_1595	m1595	(input_data_all[1796:0],output_data_all[1595]);
module_output_bit_1596	m1596	(input_data_all[1796:0],output_data_all[1596]);
module_output_bit_1597	m1597	(input_data_all[1796:0],output_data_all[1597]);
module_output_bit_1598	m1598	(input_data_all[1796:0],output_data_all[1598]);
module_output_bit_1599	m1599	(input_data_all[1796:0],output_data_all[1599]);
module_output_bit_1600	m1600	(input_data_all[1796:0],output_data_all[1600]);
module_output_bit_1601	m1601	(input_data_all[1796:0],output_data_all[1601]);
module_output_bit_1602	m1602	(input_data_all[1796:0],output_data_all[1602]);
module_output_bit_1603	m1603	(input_data_all[1796:0],output_data_all[1603]);
module_output_bit_1604	m1604	(input_data_all[1796:0],output_data_all[1604]);
module_output_bit_1605	m1605	(input_data_all[1796:0],output_data_all[1605]);
module_output_bit_1606	m1606	(input_data_all[1796:0],output_data_all[1606]);
module_output_bit_1607	m1607	(input_data_all[1796:0],output_data_all[1607]);
module_output_bit_1608	m1608	(input_data_all[1796:0],output_data_all[1608]);
module_output_bit_1609	m1609	(input_data_all[1796:0],output_data_all[1609]);
module_output_bit_1610	m1610	(input_data_all[1796:0],output_data_all[1610]);
module_output_bit_1611	m1611	(input_data_all[1796:0],output_data_all[1611]);
module_output_bit_1612	m1612	(input_data_all[1796:0],output_data_all[1612]);
module_output_bit_1613	m1613	(input_data_all[1796:0],output_data_all[1613]);
module_output_bit_1614	m1614	(input_data_all[1796:0],output_data_all[1614]);
module_output_bit_1615	m1615	(input_data_all[1796:0],output_data_all[1615]);
module_output_bit_1616	m1616	(input_data_all[1796:0],output_data_all[1616]);
module_output_bit_1617	m1617	(input_data_all[1796:0],output_data_all[1617]);
module_output_bit_1618	m1618	(input_data_all[1796:0],output_data_all[1618]);
module_output_bit_1619	m1619	(input_data_all[1796:0],output_data_all[1619]);
module_output_bit_1620	m1620	(input_data_all[1796:0],output_data_all[1620]);
module_output_bit_1621	m1621	(input_data_all[1796:0],output_data_all[1621]);
module_output_bit_1622	m1622	(input_data_all[1796:0],output_data_all[1622]);
module_output_bit_1623	m1623	(input_data_all[1796:0],output_data_all[1623]);
module_output_bit_1624	m1624	(input_data_all[1796:0],output_data_all[1624]);
module_output_bit_1625	m1625	(input_data_all[1796:0],output_data_all[1625]);
module_output_bit_1626	m1626	(input_data_all[1796:0],output_data_all[1626]);
module_output_bit_1627	m1627	(input_data_all[1796:0],output_data_all[1627]);
module_output_bit_1628	m1628	(input_data_all[1796:0],output_data_all[1628]);
module_output_bit_1629	m1629	(input_data_all[1796:0],output_data_all[1629]);
module_output_bit_1630	m1630	(input_data_all[1796:0],output_data_all[1630]);
module_output_bit_1631	m1631	(input_data_all[1796:0],output_data_all[1631]);
module_output_bit_1632	m1632	(input_data_all[1796:0],output_data_all[1632]);
module_output_bit_1633	m1633	(input_data_all[1796:0],output_data_all[1633]);
module_output_bit_1634	m1634	(input_data_all[1796:0],output_data_all[1634]);
module_output_bit_1635	m1635	(input_data_all[1796:0],output_data_all[1635]);
module_output_bit_1636	m1636	(input_data_all[1796:0],output_data_all[1636]);
module_output_bit_1637	m1637	(input_data_all[1796:0],output_data_all[1637]);
module_output_bit_1638	m1638	(input_data_all[1796:0],output_data_all[1638]);
module_output_bit_1639	m1639	(input_data_all[1796:0],output_data_all[1639]);
module_output_bit_1640	m1640	(input_data_all[1796:0],output_data_all[1640]);
module_output_bit_1641	m1641	(input_data_all[1796:0],output_data_all[1641]);
module_output_bit_1642	m1642	(input_data_all[1796:0],output_data_all[1642]);
module_output_bit_1643	m1643	(input_data_all[1796:0],output_data_all[1643]);
module_output_bit_1644	m1644	(input_data_all[1796:0],output_data_all[1644]);
module_output_bit_1645	m1645	(input_data_all[1796:0],output_data_all[1645]);
module_output_bit_1646	m1646	(input_data_all[1796:0],output_data_all[1646]);
module_output_bit_1647	m1647	(input_data_all[1796:0],output_data_all[1647]);
module_output_bit_1648	m1648	(input_data_all[1796:0],output_data_all[1648]);
module_output_bit_1649	m1649	(input_data_all[1796:0],output_data_all[1649]);
module_output_bit_1650	m1650	(input_data_all[1796:0],output_data_all[1650]);
module_output_bit_1651	m1651	(input_data_all[1796:0],output_data_all[1651]);
module_output_bit_1652	m1652	(input_data_all[1796:0],output_data_all[1652]);
module_output_bit_1653	m1653	(input_data_all[1796:0],output_data_all[1653]);
module_output_bit_1654	m1654	(input_data_all[1796:0],output_data_all[1654]);
module_output_bit_1655	m1655	(input_data_all[1796:0],output_data_all[1655]);
module_output_bit_1656	m1656	(input_data_all[1796:0],output_data_all[1656]);
module_output_bit_1657	m1657	(input_data_all[1796:0],output_data_all[1657]);
module_output_bit_1658	m1658	(input_data_all[1796:0],output_data_all[1658]);
module_output_bit_1659	m1659	(input_data_all[1796:0],output_data_all[1659]);
module_output_bit_1660	m1660	(input_data_all[1796:0],output_data_all[1660]);
module_output_bit_1661	m1661	(input_data_all[1796:0],output_data_all[1661]);
module_output_bit_1662	m1662	(input_data_all[1796:0],output_data_all[1662]);
module_output_bit_1663	m1663	(input_data_all[1796:0],output_data_all[1663]);
module_output_bit_1664	m1664	(input_data_all[1796:0],output_data_all[1664]);
module_output_bit_1665	m1665	(input_data_all[1796:0],output_data_all[1665]);
module_output_bit_1666	m1666	(input_data_all[1796:0],output_data_all[1666]);
module_output_bit_1667	m1667	(input_data_all[1796:0],output_data_all[1667]);
module_output_bit_1668	m1668	(input_data_all[1796:0],output_data_all[1668]);
module_output_bit_1669	m1669	(input_data_all[1796:0],output_data_all[1669]);
module_output_bit_1670	m1670	(input_data_all[1796:0],output_data_all[1670]);
module_output_bit_1671	m1671	(input_data_all[1796:0],output_data_all[1671]);
module_output_bit_1672	m1672	(input_data_all[1796:0],output_data_all[1672]);
module_output_bit_1673	m1673	(input_data_all[1796:0],output_data_all[1673]);
module_output_bit_1674	m1674	(input_data_all[1796:0],output_data_all[1674]);
module_output_bit_1675	m1675	(input_data_all[1796:0],output_data_all[1675]);
module_output_bit_1676	m1676	(input_data_all[1796:0],output_data_all[1676]);
module_output_bit_1677	m1677	(input_data_all[1796:0],output_data_all[1677]);
module_output_bit_1678	m1678	(input_data_all[1796:0],output_data_all[1678]);
module_output_bit_1679	m1679	(input_data_all[1796:0],output_data_all[1679]);
module_output_bit_1680	m1680	(input_data_all[1796:0],output_data_all[1680]);
module_output_bit_1681	m1681	(input_data_all[1796:0],output_data_all[1681]);
module_output_bit_1682	m1682	(input_data_all[1796:0],output_data_all[1682]);
module_output_bit_1683	m1683	(input_data_all[1796:0],output_data_all[1683]);
module_output_bit_1684	m1684	(input_data_all[1796:0],output_data_all[1684]);
module_output_bit_1685	m1685	(input_data_all[1796:0],output_data_all[1685]);
module_output_bit_1686	m1686	(input_data_all[1796:0],output_data_all[1686]);
module_output_bit_1687	m1687	(input_data_all[1796:0],output_data_all[1687]);
module_output_bit_1688	m1688	(input_data_all[1796:0],output_data_all[1688]);
module_output_bit_1689	m1689	(input_data_all[1796:0],output_data_all[1689]);
module_output_bit_1690	m1690	(input_data_all[1796:0],output_data_all[1690]);
module_output_bit_1691	m1691	(input_data_all[1796:0],output_data_all[1691]);
module_output_bit_1692	m1692	(input_data_all[1796:0],output_data_all[1692]);
module_output_bit_1693	m1693	(input_data_all[1796:0],output_data_all[1693]);
module_output_bit_1694	m1694	(input_data_all[1796:0],output_data_all[1694]);
module_output_bit_1695	m1695	(input_data_all[1796:0],output_data_all[1695]);
module_output_bit_1696	m1696	(input_data_all[1796:0],output_data_all[1696]);
module_output_bit_1697	m1697	(input_data_all[1796:0],output_data_all[1697]);
module_output_bit_1698	m1698	(input_data_all[1796:0],output_data_all[1698]);
module_output_bit_1699	m1699	(input_data_all[1796:0],output_data_all[1699]);
module_output_bit_1700	m1700	(input_data_all[1796:0],output_data_all[1700]);
module_output_bit_1701	m1701	(input_data_all[1796:0],output_data_all[1701]);
module_output_bit_1702	m1702	(input_data_all[1796:0],output_data_all[1702]);
module_output_bit_1703	m1703	(input_data_all[1796:0],output_data_all[1703]);
module_output_bit_1704	m1704	(input_data_all[1796:0],output_data_all[1704]);
module_output_bit_1705	m1705	(input_data_all[1796:0],output_data_all[1705]);
module_output_bit_1706	m1706	(input_data_all[1796:0],output_data_all[1706]);
module_output_bit_1707	m1707	(input_data_all[1796:0],output_data_all[1707]);
module_output_bit_1708	m1708	(input_data_all[1796:0],output_data_all[1708]);
module_output_bit_1709	m1709	(input_data_all[1796:0],output_data_all[1709]);
module_output_bit_1710	m1710	(input_data_all[1796:0],output_data_all[1710]);
module_output_bit_1711	m1711	(input_data_all[1796:0],output_data_all[1711]);
module_output_bit_1712	m1712	(input_data_all[1796:0],output_data_all[1712]);
module_output_bit_1713	m1713	(input_data_all[1796:0],output_data_all[1713]);
module_output_bit_1714	m1714	(input_data_all[1796:0],output_data_all[1714]);
module_output_bit_1715	m1715	(input_data_all[1796:0],output_data_all[1715]);
module_output_bit_1716	m1716	(input_data_all[1796:0],output_data_all[1716]);
module_output_bit_1717	m1717	(input_data_all[1796:0],output_data_all[1717]);
module_output_bit_1718	m1718	(input_data_all[1796:0],output_data_all[1718]);
module_output_bit_1719	m1719	(input_data_all[1796:0],output_data_all[1719]);
module_output_bit_1720	m1720	(input_data_all[1796:0],output_data_all[1720]);
module_output_bit_1721	m1721	(input_data_all[1796:0],output_data_all[1721]);
module_output_bit_1722	m1722	(input_data_all[1796:0],output_data_all[1722]);
module_output_bit_1723	m1723	(input_data_all[1796:0],output_data_all[1723]);
module_output_bit_1724	m1724	(input_data_all[1796:0],output_data_all[1724]);
module_output_bit_1725	m1725	(input_data_all[1796:0],output_data_all[1725]);
module_output_bit_1726	m1726	(input_data_all[1796:0],output_data_all[1726]);
module_output_bit_1727	m1727	(input_data_all[1796:0],output_data_all[1727]);
module_output_bit_1728	m1728	(input_data_all[1796:0],output_data_all[1728]);
module_output_bit_1729	m1729	(input_data_all[1796:0],output_data_all[1729]);
module_output_bit_1730	m1730	(input_data_all[1796:0],output_data_all[1730]);
module_output_bit_1731	m1731	(input_data_all[1796:0],output_data_all[1731]);
module_output_bit_1732	m1732	(input_data_all[1796:0],output_data_all[1732]);
module_output_bit_1733	m1733	(input_data_all[1796:0],output_data_all[1733]);
module_output_bit_1734	m1734	(input_data_all[1796:0],output_data_all[1734]);
module_output_bit_1735	m1735	(input_data_all[1796:0],output_data_all[1735]);
module_output_bit_1736	m1736	(input_data_all[1796:0],output_data_all[1736]);
module_output_bit_1737	m1737	(input_data_all[1796:0],output_data_all[1737]);
module_output_bit_1738	m1738	(input_data_all[1796:0],output_data_all[1738]);
module_output_bit_1739	m1739	(input_data_all[1796:0],output_data_all[1739]);
module_output_bit_1740	m1740	(input_data_all[1796:0],output_data_all[1740]);
module_output_bit_1741	m1741	(input_data_all[1796:0],output_data_all[1741]);
module_output_bit_1742	m1742	(input_data_all[1796:0],output_data_all[1742]);
module_output_bit_1743	m1743	(input_data_all[1796:0],output_data_all[1743]);
module_output_bit_1744	m1744	(input_data_all[1796:0],output_data_all[1744]);
module_output_bit_1745	m1745	(input_data_all[1796:0],output_data_all[1745]);
module_output_bit_1746	m1746	(input_data_all[1796:0],output_data_all[1746]);
module_output_bit_1747	m1747	(input_data_all[1796:0],output_data_all[1747]);
module_output_bit_1748	m1748	(input_data_all[1796:0],output_data_all[1748]);
module_output_bit_1749	m1749	(input_data_all[1796:0],output_data_all[1749]);
module_output_bit_1750	m1750	(input_data_all[1796:0],output_data_all[1750]);
module_output_bit_1751	m1751	(input_data_all[1796:0],output_data_all[1751]);
module_output_bit_1752	m1752	(input_data_all[1796:0],output_data_all[1752]);
module_output_bit_1753	m1753	(input_data_all[1796:0],output_data_all[1753]);
module_output_bit_1754	m1754	(input_data_all[1796:0],output_data_all[1754]);
module_output_bit_1755	m1755	(input_data_all[1796:0],output_data_all[1755]);
module_output_bit_1756	m1756	(input_data_all[1796:0],output_data_all[1756]);
module_output_bit_1757	m1757	(input_data_all[1796:0],output_data_all[1757]);
module_output_bit_1758	m1758	(input_data_all[1796:0],output_data_all[1758]);
module_output_bit_1759	m1759	(input_data_all[1796:0],output_data_all[1759]);
module_output_bit_1760	m1760	(input_data_all[1796:0],output_data_all[1760]);
module_output_bit_1761	m1761	(input_data_all[1796:0],output_data_all[1761]);
module_output_bit_1762	m1762	(input_data_all[1796:0],output_data_all[1762]);
module_output_bit_1763	m1763	(input_data_all[1796:0],output_data_all[1763]);
module_output_bit_1764	m1764	(input_data_all[1796:0],output_data_all[1764]);
module_output_bit_1765	m1765	(input_data_all[1796:0],output_data_all[1765]);
module_output_bit_1766	m1766	(input_data_all[1796:0],output_data_all[1766]);
module_output_bit_1767	m1767	(input_data_all[1796:0],output_data_all[1767]);
module_output_bit_1768	m1768	(input_data_all[1796:0],output_data_all[1768]);
module_output_bit_1769	m1769	(input_data_all[1796:0],output_data_all[1769]);
module_output_bit_1770	m1770	(input_data_all[1796:0],output_data_all[1770]);
module_output_bit_1771	m1771	(input_data_all[1796:0],output_data_all[1771]);
module_output_bit_1772	m1772	(input_data_all[1796:0],output_data_all[1772]);
module_output_bit_1773	m1773	(input_data_all[1796:0],output_data_all[1773]);
module_output_bit_1774	m1774	(input_data_all[1796:0],output_data_all[1774]);
module_output_bit_1775	m1775	(input_data_all[1796:0],output_data_all[1775]);
module_output_bit_1776	m1776	(input_data_all[1796:0],output_data_all[1776]);
module_output_bit_1777	m1777	(input_data_all[1796:0],output_data_all[1777]);
module_output_bit_1778	m1778	(input_data_all[1796:0],output_data_all[1778]);
module_output_bit_1779	m1779	(input_data_all[1796:0],output_data_all[1779]);
module_output_bit_1780	m1780	(input_data_all[1796:0],output_data_all[1780]);
module_output_bit_1781	m1781	(input_data_all[1796:0],output_data_all[1781]);
module_output_bit_1782	m1782	(input_data_all[1796:0],output_data_all[1782]);
module_output_bit_1783	m1783	(input_data_all[1796:0],output_data_all[1783]);
module_output_bit_1784	m1784	(input_data_all[1796:0],output_data_all[1784]);
module_output_bit_1785	m1785	(input_data_all[1796:0],output_data_all[1785]);
module_output_bit_1786	m1786	(input_data_all[1796:0],output_data_all[1786]);
module_output_bit_1787	m1787	(input_data_all[1796:0],output_data_all[1787]);
module_output_bit_1788	m1788	(input_data_all[1796:0],output_data_all[1788]);
module_output_bit_1789	m1789	(input_data_all[1796:0],output_data_all[1789]);
module_output_bit_1790	m1790	(input_data_all[1796:0],output_data_all[1790]);
module_output_bit_1791	m1791	(input_data_all[1796:0],output_data_all[1791]);
module_output_bit_1792	m1792	(input_data_all[1796:0],output_data_all[1792]);
module_output_bit_1793	m1793	(input_data_all[1796:0],output_data_all[1793]);
module_output_bit_1794	m1794	(input_data_all[1796:0],output_data_all[1794]);
module_output_bit_1795	m1795	(input_data_all[1796:0],output_data_all[1795]);
module_output_bit_1796	m1796	(input_data_all[1796:0],output_data_all[1796]);
module_output_bit_1797	m1797	(input_data_all[1796:0],output_data_all[1797]);
module_output_bit_1798	m1798	(input_data_all[1796:0],output_data_all[1798]);
module_output_bit_1799	m1799	(input_data_all[1796:0],output_data_all[1799]);
module_output_bit_1800	m1800	(input_data_all[1796:0],output_data_all[1800]);
module_output_bit_1801	m1801	(input_data_all[1796:0],output_data_all[1801]);
module_output_bit_1802	m1802	(input_data_all[1796:0],output_data_all[1802]);
module_output_bit_1803	m1803	(input_data_all[1796:0],output_data_all[1803]);
module_output_bit_1804	m1804	(input_data_all[1796:0],output_data_all[1804]);
module_output_bit_1805	m1805	(input_data_all[1796:0],output_data_all[1805]);
module_output_bit_1806	m1806	(input_data_all[1796:0],output_data_all[1806]);
module_output_bit_1807	m1807	(input_data_all[1796:0],output_data_all[1807]);
module_output_bit_1808	m1808	(input_data_all[1796:0],output_data_all[1808]);
module_output_bit_1809	m1809	(input_data_all[1796:0],output_data_all[1809]);
module_output_bit_1810	m1810	(input_data_all[1796:0],output_data_all[1810]);
module_output_bit_1811	m1811	(input_data_all[1796:0],output_data_all[1811]);
module_output_bit_1812	m1812	(input_data_all[1796:0],output_data_all[1812]);
module_output_bit_1813	m1813	(input_data_all[1796:0],output_data_all[1813]);
module_output_bit_1814	m1814	(input_data_all[1796:0],output_data_all[1814]);
module_output_bit_1815	m1815	(input_data_all[1796:0],output_data_all[1815]);
module_output_bit_1816	m1816	(input_data_all[1796:0],output_data_all[1816]);
module_output_bit_1817	m1817	(input_data_all[1796:0],output_data_all[1817]);
module_output_bit_1818	m1818	(input_data_all[1796:0],output_data_all[1818]);
module_output_bit_1819	m1819	(input_data_all[1796:0],output_data_all[1819]);
module_output_bit_1820	m1820	(input_data_all[1796:0],output_data_all[1820]);
module_output_bit_1821	m1821	(input_data_all[1796:0],output_data_all[1821]);
module_output_bit_1822	m1822	(input_data_all[1796:0],output_data_all[1822]);
module_output_bit_1823	m1823	(input_data_all[1796:0],output_data_all[1823]);
module_output_bit_1824	m1824	(input_data_all[1796:0],output_data_all[1824]);
module_output_bit_1825	m1825	(input_data_all[1796:0],output_data_all[1825]);

endmodule