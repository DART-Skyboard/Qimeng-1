//circuit accuracy = 1
//test amounts  = 1000000
//total BDD nodes = 33224
//total split modes = 20587
//train time = 9408.04
module module_output_bit_63(i,o);

input [1893:0] i;
output  o;

wire [0:0] l_0;
wire [1:0] l_1;
wire [3:0] l_2;
wire [7:0] l_3;
wire [13:0] l_4;
wire [13:0] l_5;
wire [13:0] l_6;
wire [13:0] l_7;
wire [19:0] l_8;
wire [17:0] l_9;
wire [17:0] l_10;
wire [17:0] l_11;
wire [17:0] l_12;
wire [17:0] l_13;
wire [17:0] l_14;
wire [17:0] l_15;
wire [17:0] l_16;
wire [12:0] l_17;
wire [12:0] l_18;
wire [18:0] l_19;
wire [23:0] l_20;
wire [23:0] l_21;
wire [27:0] l_22;
wire [35:0] l_23;
wire [51:0] l_24;
wire [53:0] l_25;
wire [85:0] l_26;
wire [89:0] l_27;
wire [97:0] l_28;
wire [113:0] l_29;
wire [145:0] l_30;
wire [209:0] l_31;
wire [273:0] l_32;
wire [401:0] l_33;
wire [529:0] l_34;
wire [785:0] l_35;
wire [1041:0] l_36;
wire [1553:0] l_37;
wire [2065:0] l_38;
wire [3089:0] l_39;
wire [4113:0] l_40;
wire [6177:0] l_41;
wire [8257:0] l_42;
wire [414:0] l_43;
wire [281:0] l_44;
wire [393:0] l_45;
wire [536:0] l_46;
wire [1063:0] l_47;
wire [548:0] l_48;
wire [141:0] l_49;
wire [76:0] l_50;
wire [43:0] l_51;
wire [74:0] l_52;
wire [41:0] l_53;
wire [24:0] l_54;
wire [15:0] l_55;
wire [14:0] l_56;
wire [6:0] l_57;
wire [2:0] l_58;
wire [0:0] l_59;
wire [-1:0] l_60;

assign o = l_0[0];

assign l_0[0]    = ( l_1 [0] & !i[63]) | ( l_1 [1] &  i[63]);
assign l_1[0]    = ( l_2 [0] & !i[1713]) | ( l_2 [1] &  i[1713]);
assign l_1[1]    = ( l_2 [2] & !i[1713]) | ( l_2 [3] &  i[1713]);
assign l_2[0]    = ( l_3 [0] & !i[1714]) | ( l_3 [1] &  i[1714]);
assign l_2[1]    = ( l_3 [2] & !i[1714]) | ( l_3 [3] &  i[1714]);
assign l_2[2]    = ( l_3 [4] & !i[1714]) | ( l_3 [5] &  i[1714]);
assign l_2[3]    = ( l_3 [6] & !i[1714]) | ( l_3 [7] &  i[1714]);
assign l_3[0]    = ( l_4 [0] &  i[1715]);
assign l_3[1]    = ( l_4 [1] & !i[1715]) | ( l_4 [2] &  i[1715]);
assign l_3[2]    = ( l_4 [3] & !i[1715]) | ( l_4 [4] &  i[1715]);
assign l_3[3]    = ( l_4 [5] & !i[1715]) | ( l_4 [6] &  i[1715]);
assign l_3[4]    = (!i[1715]) | ( l_4 [7] &  i[1715]);
assign l_3[5]    = ( l_4 [8] & !i[1715]) | ( l_4 [9] &  i[1715]);
assign l_3[6]    = ( l_4 [10] & !i[1715]) | ( l_4 [11] &  i[1715]);
assign l_3[7]    = ( l_4 [12] & !i[1715]) | ( l_4 [13] &  i[1715]);
assign l_4[0]    = ( l_5 [0] & !i[1716]);
assign l_4[1]    = ( l_5 [1] & !i[1716]);
assign l_4[2]    = ( l_5 [2] & !i[1716]);
assign l_4[3]    = ( l_5 [3] & !i[1716]);
assign l_4[4]    = ( l_5 [4] & !i[1716]);
assign l_4[5]    = ( l_5 [5] & !i[1716]);
assign l_4[6]    = ( l_5 [6] & !i[1716]);
assign l_4[7]    = ( l_5 [7] & !i[1716]) | (      i[1716]);
assign l_4[8]    = ( l_5 [8] & !i[1716]) | (      i[1716]);
assign l_4[9]    = ( l_5 [9] & !i[1716]) | (      i[1716]);
assign l_4[10]    = ( l_5 [10] & !i[1716]) | (      i[1716]);
assign l_4[11]    = ( l_5 [11] & !i[1716]) | (      i[1716]);
assign l_4[12]    = ( l_5 [12] & !i[1716]) | (      i[1716]);
assign l_4[13]    = ( l_5 [13] & !i[1716]) | (      i[1716]);
assign l_5[0]    = ( l_6 [0] & !i[1717]);
assign l_5[1]    = ( l_6 [1] & !i[1717]);
assign l_5[2]    = ( l_6 [2] & !i[1717]);
assign l_5[3]    = ( l_6 [3] & !i[1717]);
assign l_5[4]    = ( l_6 [4] & !i[1717]);
assign l_5[5]    = ( l_6 [5] & !i[1717]);
assign l_5[6]    = ( l_6 [6] & !i[1717]);
assign l_5[7]    = ( l_6 [7] & !i[1717]) | (      i[1717]);
assign l_5[8]    = ( l_6 [8] & !i[1717]) | (      i[1717]);
assign l_5[9]    = ( l_6 [9] & !i[1717]) | (      i[1717]);
assign l_5[10]    = ( l_6 [10] & !i[1717]) | (      i[1717]);
assign l_5[11]    = ( l_6 [11] & !i[1717]) | (      i[1717]);
assign l_5[12]    = ( l_6 [12] & !i[1717]) | (      i[1717]);
assign l_5[13]    = ( l_6 [13] & !i[1717]) | (      i[1717]);
assign l_6[0]    = ( l_7 [0] &  i[1723]);
assign l_6[1]    = ( l_7 [1] &  i[1723]);
assign l_6[2]    = ( l_7 [2] &  i[1723]);
assign l_6[3]    = ( l_7 [3] &  i[1723]);
assign l_6[4]    = ( l_7 [4] &  i[1723]);
assign l_6[5]    = ( l_7 [5] &  i[1723]);
assign l_6[6]    = ( l_7 [6] &  i[1723]);
assign l_6[7]    = (!i[1723]) | ( l_7 [7] &  i[1723]);
assign l_6[8]    = (!i[1723]) | ( l_7 [8] &  i[1723]);
assign l_6[9]    = (!i[1723]) | ( l_7 [9] &  i[1723]);
assign l_6[10]    = (!i[1723]) | ( l_7 [10] &  i[1723]);
assign l_6[11]    = (!i[1723]) | ( l_7 [11] &  i[1723]);
assign l_6[12]    = (!i[1723]) | ( l_7 [12] &  i[1723]);
assign l_6[13]    = (!i[1723]) | ( l_7 [13] &  i[1723]);
assign l_7[0]    = ( l_8 [0] & !i[1707]);
assign l_7[1]    = ( l_8 [1] & !i[1707]) | ( l_8 [2] &  i[1707]);
assign l_7[2]    = ( l_8 [3] & !i[1707]) | ( l_8 [4] &  i[1707]);
assign l_7[3]    = ( l_8 [5] & !i[1707]) | ( l_8 [6] &  i[1707]);
assign l_7[4]    = ( l_8 [7] & !i[1707]) | ( l_8 [8] &  i[1707]);
assign l_7[5]    = ( l_8 [5] & !i[1707]) | ( l_8 [9] &  i[1707]);
assign l_7[6]    = ( l_8 [5] &  i[1707]);
assign l_7[7]    = ( l_8 [10] & !i[1707]) | ( l_8 [11] &  i[1707]);
assign l_7[8]    = ( l_8 [12] & !i[1707]) | ( l_8 [13] &  i[1707]);
assign l_7[9]    = ( l_8 [14] & !i[1707]) | ( l_8 [15] &  i[1707]);
assign l_7[10]    = (!l_8 [6] & !i[1707]) | ( l_8 [16] &  i[1707]);
assign l_7[11]    = ( l_8 [17] & !i[1707]) | ( l_8 [18] &  i[1707]);
assign l_7[12]    = (!l_8 [6] & !i[1707]) | (      i[1707]);
assign l_7[13]    = (!l_8 [9] & !i[1707]) | ( l_8 [19] &  i[1707]);
assign l_8[0]    = ( l_9 [0] & !i[1724]);
assign l_8[1]    = ( l_9 [1] & !i[1724]);
assign l_8[2]    = ( l_9 [2] & !i[1724]);
assign l_8[3]    = ( l_9 [3] & !i[1724]);
assign l_8[4]    = ( l_9 [4] & !i[1724]);
assign l_8[5]    = ( l_9 [5] & !i[1724]);
assign l_8[6]    = ( l_9 [6] & !i[1724]);
assign l_8[7]    = ( l_9 [7] & !i[1724]);
assign l_8[8]    = ( l_9 [8] & !i[1724]);
assign l_8[9]    = ( l_9 [9] & !i[1724]);
assign l_8[10]    = ( l_9 [10] & !i[1724]) | (      i[1724]);
assign l_8[11]    = ( l_9 [11] & !i[1724]) | (      i[1724]);
assign l_8[12]    = ( l_9 [12] & !i[1724]) | (      i[1724]);
assign l_8[13]    = ( l_9 [13] & !i[1724]) | (      i[1724]);
assign l_8[14]    = ( l_9 [14] & !i[1724]) | (      i[1724]);
assign l_8[15]    = ( l_9 [15] & !i[1724]) | (      i[1724]);
assign l_8[16]    = (!l_9 [5] & !i[1724]) | (      i[1724]);
assign l_8[17]    = ( l_9 [16] & !i[1724]) | (      i[1724]);
assign l_8[18]    = ( l_9 [17] & !i[1724]) | (      i[1724]);
assign l_8[19]    = (!l_9 [6] & !i[1724]) | (      i[1724]);
assign l_9[0]    = ( l_10 [0] & !i[1721]);
assign l_9[1]    = ( l_10 [1] & !i[1721]);
assign l_9[2]    = ( l_10 [2] & !i[1721]);
assign l_9[3]    = ( l_10 [3] & !i[1721]);
assign l_9[4]    = ( l_10 [4] & !i[1721]);
assign l_9[5]    = ( l_10 [5] & !i[1721]);
assign l_9[6]    = ( l_10 [6] & !i[1721]);
assign l_9[7]    = ( l_10 [7] & !i[1721]);
assign l_9[8]    = ( l_10 [8] & !i[1721]);
assign l_9[9]    = ( l_10 [9] & !i[1721]);
assign l_9[10]    = ( l_10 [10] & !i[1721]) | (      i[1721]);
assign l_9[11]    = ( l_10 [11] & !i[1721]) | (      i[1721]);
assign l_9[12]    = ( l_10 [12] & !i[1721]) | (      i[1721]);
assign l_9[13]    = ( l_10 [13] & !i[1721]) | (      i[1721]);
assign l_9[14]    = ( l_10 [14] & !i[1721]) | (      i[1721]);
assign l_9[15]    = ( l_10 [15] & !i[1721]) | (      i[1721]);
assign l_9[16]    = ( l_10 [16] & !i[1721]) | (      i[1721]);
assign l_9[17]    = ( l_10 [17] & !i[1721]) | (      i[1721]);
assign l_10[0]    = ( l_11 [0] &  i[1726]);
assign l_10[1]    = ( l_11 [1] &  i[1726]);
assign l_10[2]    = ( l_11 [2] &  i[1726]);
assign l_10[3]    = ( l_11 [3] &  i[1726]);
assign l_10[4]    = ( l_11 [4] &  i[1726]);
assign l_10[5]    = ( l_11 [5] &  i[1726]);
assign l_10[6]    = ( l_11 [6] &  i[1726]);
assign l_10[7]    = ( l_11 [7] &  i[1726]);
assign l_10[8]    = ( l_11 [8] &  i[1726]);
assign l_10[9]    = ( l_11 [9] &  i[1726]);
assign l_10[10]    = (!i[1726]) | ( l_11 [10] &  i[1726]);
assign l_10[11]    = (!i[1726]) | ( l_11 [11] &  i[1726]);
assign l_10[12]    = (!i[1726]) | ( l_11 [12] &  i[1726]);
assign l_10[13]    = (!i[1726]) | ( l_11 [13] &  i[1726]);
assign l_10[14]    = (!i[1726]) | ( l_11 [14] &  i[1726]);
assign l_10[15]    = (!i[1726]) | ( l_11 [15] &  i[1726]);
assign l_10[16]    = (!i[1726]) | ( l_11 [16] &  i[1726]);
assign l_10[17]    = (!i[1726]) | ( l_11 [17] &  i[1726]);
assign l_11[0]    = ( l_12 [0] &  i[1727]);
assign l_11[1]    = ( l_12 [1] &  i[1727]);
assign l_11[2]    = ( l_12 [2] &  i[1727]);
assign l_11[3]    = ( l_12 [3] &  i[1727]);
assign l_11[4]    = ( l_12 [4] &  i[1727]);
assign l_11[5]    = ( l_12 [5] &  i[1727]);
assign l_11[6]    = ( l_12 [6] &  i[1727]);
assign l_11[7]    = ( l_12 [7] &  i[1727]);
assign l_11[8]    = ( l_12 [8] &  i[1727]);
assign l_11[9]    = ( l_12 [9] &  i[1727]);
assign l_11[10]    = (!i[1727]) | ( l_12 [10] &  i[1727]);
assign l_11[11]    = (!i[1727]) | ( l_12 [11] &  i[1727]);
assign l_11[12]    = (!i[1727]) | ( l_12 [12] &  i[1727]);
assign l_11[13]    = (!i[1727]) | ( l_12 [13] &  i[1727]);
assign l_11[14]    = (!i[1727]) | ( l_12 [14] &  i[1727]);
assign l_11[15]    = (!i[1727]) | ( l_12 [15] &  i[1727]);
assign l_11[16]    = (!i[1727]) | ( l_12 [16] &  i[1727]);
assign l_11[17]    = (!i[1727]) | ( l_12 [17] &  i[1727]);
assign l_12[0]    = ( l_13 [0] & !i[1725]);
assign l_12[1]    = ( l_13 [1] & !i[1725]);
assign l_12[2]    = ( l_13 [2] & !i[1725]);
assign l_12[3]    = ( l_13 [3] & !i[1725]);
assign l_12[4]    = ( l_13 [4] & !i[1725]);
assign l_12[5]    = ( l_13 [5] & !i[1725]);
assign l_12[6]    = ( l_13 [6] & !i[1725]);
assign l_12[7]    = ( l_13 [7] & !i[1725]);
assign l_12[8]    = ( l_13 [8] & !i[1725]);
assign l_12[9]    = ( l_13 [9] & !i[1725]);
assign l_12[10]    = ( l_13 [10] & !i[1725]) | (      i[1725]);
assign l_12[11]    = ( l_13 [11] & !i[1725]) | (      i[1725]);
assign l_12[12]    = ( l_13 [12] & !i[1725]) | (      i[1725]);
assign l_12[13]    = ( l_13 [13] & !i[1725]) | (      i[1725]);
assign l_12[14]    = ( l_13 [14] & !i[1725]) | (      i[1725]);
assign l_12[15]    = ( l_13 [15] & !i[1725]) | (      i[1725]);
assign l_12[16]    = ( l_13 [16] & !i[1725]) | (      i[1725]);
assign l_12[17]    = ( l_13 [17] & !i[1725]) | (      i[1725]);
assign l_13[0]    = ( l_14 [0] & !i[1722]);
assign l_13[1]    = ( l_14 [1] & !i[1722]);
assign l_13[2]    = ( l_14 [2] & !i[1722]);
assign l_13[3]    = ( l_14 [3] & !i[1722]);
assign l_13[4]    = ( l_14 [4] & !i[1722]);
assign l_13[5]    = ( l_14 [5] & !i[1722]);
assign l_13[6]    = ( l_14 [6] & !i[1722]);
assign l_13[7]    = ( l_14 [7] & !i[1722]);
assign l_13[8]    = ( l_14 [8] & !i[1722]);
assign l_13[9]    = ( l_14 [9] & !i[1722]);
assign l_13[10]    = ( l_14 [10] & !i[1722]) | (      i[1722]);
assign l_13[11]    = ( l_14 [11] & !i[1722]) | (      i[1722]);
assign l_13[12]    = ( l_14 [12] & !i[1722]) | (      i[1722]);
assign l_13[13]    = ( l_14 [13] & !i[1722]) | (      i[1722]);
assign l_13[14]    = ( l_14 [14] & !i[1722]) | (      i[1722]);
assign l_13[15]    = ( l_14 [15] & !i[1722]) | (      i[1722]);
assign l_13[16]    = ( l_14 [16] & !i[1722]) | (      i[1722]);
assign l_13[17]    = ( l_14 [17] & !i[1722]) | (      i[1722]);
assign l_14[0]    = ( l_15 [0] & !i[1718]);
assign l_14[1]    = ( l_15 [1] & !i[1718]);
assign l_14[2]    = ( l_15 [2] & !i[1718]);
assign l_14[3]    = ( l_15 [3] & !i[1718]);
assign l_14[4]    = ( l_15 [4] & !i[1718]);
assign l_14[5]    = ( l_15 [5] & !i[1718]);
assign l_14[6]    = ( l_15 [6] & !i[1718]);
assign l_14[7]    = ( l_15 [7] & !i[1718]);
assign l_14[8]    = ( l_15 [8] & !i[1718]);
assign l_14[9]    = ( l_15 [9] & !i[1718]);
assign l_14[10]    = ( l_15 [10] & !i[1718]) | (      i[1718]);
assign l_14[11]    = ( l_15 [11] & !i[1718]) | (      i[1718]);
assign l_14[12]    = ( l_15 [12] & !i[1718]) | (      i[1718]);
assign l_14[13]    = ( l_15 [13] & !i[1718]) | (      i[1718]);
assign l_14[14]    = ( l_15 [14] & !i[1718]) | (      i[1718]);
assign l_14[15]    = ( l_15 [15] & !i[1718]) | (      i[1718]);
assign l_14[16]    = ( l_15 [16] & !i[1718]) | (      i[1718]);
assign l_14[17]    = ( l_15 [17] & !i[1718]) | (      i[1718]);
assign l_15[0]    = ( l_16 [0] & !i[1719]);
assign l_15[1]    = ( l_16 [1] & !i[1719]);
assign l_15[2]    = ( l_16 [2] & !i[1719]);
assign l_15[3]    = ( l_16 [3] & !i[1719]);
assign l_15[4]    = ( l_16 [4] & !i[1719]);
assign l_15[5]    = ( l_16 [5] & !i[1719]);
assign l_15[6]    = ( l_16 [6] & !i[1719]);
assign l_15[7]    = ( l_16 [7] & !i[1719]);
assign l_15[8]    = ( l_16 [8] & !i[1719]);
assign l_15[9]    = ( l_16 [9] & !i[1719]);
assign l_15[10]    = ( l_16 [10] & !i[1719]) | (      i[1719]);
assign l_15[11]    = ( l_16 [11] & !i[1719]) | (      i[1719]);
assign l_15[12]    = ( l_16 [12] & !i[1719]) | (      i[1719]);
assign l_15[13]    = ( l_16 [13] & !i[1719]) | (      i[1719]);
assign l_15[14]    = ( l_16 [14] & !i[1719]) | (      i[1719]);
assign l_15[15]    = ( l_16 [15] & !i[1719]) | (      i[1719]);
assign l_15[16]    = ( l_16 [16] & !i[1719]) | (      i[1719]);
assign l_15[17]    = ( l_16 [17] & !i[1719]) | (      i[1719]);
assign l_16[0]    = ( l_17 [0] &  i[1720]);
assign l_16[1]    = ( l_17 [1] &  i[1720]);
assign l_16[2]    = ( l_17 [2] &  i[1720]);
assign l_16[3]    = ( l_17 [3] &  i[1720]);
assign l_16[4]    = ( l_17 [4] &  i[1720]);
assign l_16[5]    = ( l_17 [5] &  i[1720]);
assign l_16[6]    = ( l_17 [6] &  i[1720]);
assign l_16[7]    = ( l_17 [7] &  i[1720]);
assign l_16[8]    = ( l_17 [8] &  i[1720]);
assign l_16[9]    =  i[1720];
assign l_16[10]    = (!i[1720]) | ( l_17 [9] &  i[1720]);
assign l_16[11]    = (!i[1720]) | ( l_17 [10] &  i[1720]);
assign l_16[12]    = (!i[1720]) | ( l_17 [1] &  i[1720]);
assign l_16[13]    = (!i[1720]) | ( l_17 [2] &  i[1720]);
assign l_16[14]    = (!i[1720]) | ( l_17 [3] &  i[1720]);
assign l_16[15]    = (!i[1720]) | ( l_17 [4] &  i[1720]);
assign l_16[16]    = (!i[1720]) | ( l_17 [11] &  i[1720]);
assign l_16[17]    = (!i[1720]) | ( l_17 [12] &  i[1720]);
assign l_17[0]    = ( l_18 [0] &  i[1829]);
assign l_17[1]    = ( l_18 [1]);
assign l_17[2]    = ( l_18 [2] & !i[1829]) | ( l_18 [1] &  i[1829]);
assign l_17[3]    = ( l_18 [3]);
assign l_17[4]    = ( l_18 [4] & !i[1829]) | ( l_18 [3] &  i[1829]);
assign l_17[5]    =  i[1829];
assign l_17[6]    = !i[1829];
assign l_17[7]    = ( l_18 [5] & !i[1829]) | ( l_18 [6] &  i[1829]);
assign l_17[8]    = ( l_18 [7]);
assign l_17[9]    = ( l_18 [8] & !i[1829]) | ( l_18 [9] &  i[1829]);
assign l_17[10]    = ( l_18 [8]);
assign l_17[11]    = ( l_18 [10] & !i[1829]) | ( l_18 [11] &  i[1829]);
assign l_17[12]    = ( l_18 [12]);
assign l_18[0]    = ( l_19 [0]);
assign l_18[1]    = ( l_19 [1] & !i[1798]) | ( l_19 [2] &  i[1798]);
assign l_18[2]    = ( l_19 [3] & !i[1798]) | ( l_19 [4] &  i[1798]);
assign l_18[3]    = ( l_19 [5] & !i[1798]) | ( l_19 [6] &  i[1798]);
assign l_18[4]    = ( l_19 [7] & !i[1798]) | ( l_19 [8] &  i[1798]);
assign l_18[5]    = ( l_19 [9]);
assign l_18[6]    = ( l_19 [10]);
assign l_18[7]    = ( l_19 [11] & !i[1798]) | ( l_19 [12] &  i[1798]);
assign l_18[8]    = ( l_19 [13]);
assign l_18[9]    = ( l_19 [14]);
assign l_18[10]    = ( l_19 [15]);
assign l_18[11]    = ( l_19 [16]);
assign l_18[12]    = ( l_19 [17] & !i[1798]) | ( l_19 [18] &  i[1798]);
assign l_19[0]    = ( l_20 [0]);
assign l_19[1]    = ( l_20 [1] & !i[1809]);
assign l_19[2]    = (!i[1809]) | ( l_20 [2] &  i[1809]);
assign l_19[3]    = ( l_20 [3] & !i[1809]);
assign l_19[4]    = (!i[1809]) | ( l_20 [4] &  i[1809]);
assign l_19[5]    = ( l_20 [5] & !i[1809]) | ( l_20 [6] &  i[1809]);
assign l_19[6]    = ( l_20 [6] & !i[1809]) | ( l_20 [7] &  i[1809]);
assign l_19[7]    = ( l_20 [8] & !i[1809]) | ( l_20 [6] &  i[1809]);
assign l_19[8]    = ( l_20 [6] & !i[1809]) | ( l_20 [9] &  i[1809]);
assign l_19[9]    = ( l_20 [10] & !i[1809]) | ( l_20 [11] &  i[1809]);
assign l_19[10]    = ( l_20 [12] & !i[1809]) | ( l_20 [13] &  i[1809]);
assign l_19[11]    = ( l_20 [14]);
assign l_19[12]    = ( l_20 [15]);
assign l_19[13]    = ( l_20 [16]);
assign l_19[14]    = ( l_20 [17]);
assign l_19[15]    = ( l_20 [18] & !i[1809]) | ( l_20 [19] &  i[1809]);
assign l_19[16]    = ( l_20 [20] & !i[1809]) | ( l_20 [21] &  i[1809]);
assign l_19[17]    = ( l_20 [22]);
assign l_19[18]    = ( l_20 [23]);
assign l_20[0]    = ( l_21 [0] & !i[1702]);
assign l_20[1]    = ( l_21 [1] & !i[1702]) | ( l_21 [2] &  i[1702]);
assign l_20[2]    = ( l_21 [3] & !i[1702]) | ( l_21 [4] &  i[1702]);
assign l_20[3]    = ( l_21 [5] & !i[1702]) | ( l_21 [6] &  i[1702]);
assign l_20[4]    = ( l_21 [7] & !i[1702]) | ( l_21 [8] &  i[1702]);
assign l_20[5]    = ( l_21 [9] & !i[1702]) | ( l_21 [10] &  i[1702]);
assign l_20[6]    = ( l_21 [11]);
assign l_20[7]    = ( l_21 [12] & !i[1702]) | ( l_21 [13] &  i[1702]);
assign l_20[8]    = ( l_21 [14] & !i[1702]) | ( l_21 [15] &  i[1702]);
assign l_20[9]    = ( l_21 [16] & !i[1702]) | ( l_21 [17] &  i[1702]);
assign l_20[10]    = ( l_21 [18] & !i[1702]);
assign l_20[11]    = ( l_21 [19] & !i[1702]);
assign l_20[12]    = ( l_21 [20] & !i[1702]);
assign l_20[13]    = ( l_21 [21] & !i[1702]);
assign l_20[14]    = ( l_21 [22] & !i[1702]);
assign l_20[15]    = ( l_21 [23] & !i[1702]);
assign l_20[16]    =  i[1702];
assign l_20[17]    = ( l_21 [0] & !i[1702]) | (      i[1702]);
assign l_20[18]    = ( l_21 [18] & !i[1702]) | (      i[1702]);
assign l_20[19]    = ( l_21 [19] & !i[1702]) | (      i[1702]);
assign l_20[20]    = ( l_21 [20] & !i[1702]) | (      i[1702]);
assign l_20[21]    = ( l_21 [21] & !i[1702]) | (      i[1702]);
assign l_20[22]    = ( l_21 [22] & !i[1702]) | (      i[1702]);
assign l_20[23]    = ( l_21 [23] & !i[1702]) | (      i[1702]);
assign l_21[0]    = ( l_22 [0]);
assign l_21[1]    = ( l_22 [1] & !i[1803]);
assign l_21[2]    = ( l_22 [2] & !i[1803]);
assign l_21[3]    = (!i[1803]) | ( l_22 [3] &  i[1803]);
assign l_21[4]    = (!i[1803]) | ( l_22 [4] &  i[1803]);
assign l_21[5]    = ( l_22 [5] & !i[1803]);
assign l_21[6]    = ( l_22 [6] & !i[1803]);
assign l_21[7]    = (!i[1803]) | ( l_22 [7] &  i[1803]);
assign l_21[8]    = (!i[1803]) | ( l_22 [8] &  i[1803]);
assign l_21[9]    = ( l_22 [9] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[10]    = ( l_22 [11] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[11]    = ( l_22 [10]);
assign l_21[12]    = ( l_22 [10] & !i[1803]) | ( l_22 [12] &  i[1803]);
assign l_21[13]    = ( l_22 [10] & !i[1803]) | ( l_22 [13] &  i[1803]);
assign l_21[14]    = ( l_22 [14] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[15]    = ( l_22 [15] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[16]    = ( l_22 [10] & !i[1803]) | ( l_22 [16] &  i[1803]);
assign l_21[17]    = ( l_22 [10] & !i[1803]) | ( l_22 [17] &  i[1803]);
assign l_21[18]    = ( l_22 [18] & !i[1803]) | ( l_22 [19] &  i[1803]);
assign l_21[19]    = ( l_22 [20] & !i[1803]) | ( l_22 [21] &  i[1803]);
assign l_21[20]    = ( l_22 [22] & !i[1803]) | ( l_22 [23] &  i[1803]);
assign l_21[21]    = ( l_22 [24] & !i[1803]) | ( l_22 [25] &  i[1803]);
assign l_21[22]    = ( l_22 [26]);
assign l_21[23]    = ( l_22 [27]);
assign l_22[0]    = ( l_23 [0]);
assign l_22[1]    = ( l_23 [1] & !i[1801]);
assign l_22[2]    = ( l_23 [2] & !i[1801]);
assign l_22[3]    = (!i[1801]) | ( l_23 [3] &  i[1801]);
assign l_22[4]    = (!i[1801]) | ( l_23 [4] &  i[1801]);
assign l_22[5]    = ( l_23 [5] & !i[1801]);
assign l_22[6]    = ( l_23 [6] & !i[1801]);
assign l_22[7]    = (!i[1801]) | ( l_23 [7] &  i[1801]);
assign l_22[8]    = (!i[1801]) | ( l_23 [8] &  i[1801]);
assign l_22[9]    = ( l_23 [9] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[10]    = ( l_23 [10]);
assign l_22[11]    = ( l_23 [11] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[12]    = ( l_23 [10] & !i[1801]) | ( l_23 [12] &  i[1801]);
assign l_22[13]    = ( l_23 [10] & !i[1801]) | ( l_23 [13] &  i[1801]);
assign l_22[14]    = ( l_23 [14] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[15]    = ( l_23 [15] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[16]    = ( l_23 [10] & !i[1801]) | ( l_23 [16] &  i[1801]);
assign l_22[17]    = ( l_23 [10] & !i[1801]) | ( l_23 [17] &  i[1801]);
assign l_22[18]    = ( l_23 [18] & !i[1801]) | ( l_23 [19] &  i[1801]);
assign l_22[19]    = ( l_23 [20] & !i[1801]) | ( l_23 [21] &  i[1801]);
assign l_22[20]    = ( l_23 [22] & !i[1801]) | ( l_23 [23] &  i[1801]);
assign l_22[21]    = ( l_23 [24] & !i[1801]) | ( l_23 [25] &  i[1801]);
assign l_22[22]    = ( l_23 [26] & !i[1801]) | ( l_23 [27] &  i[1801]);
assign l_22[23]    = ( l_23 [28] & !i[1801]) | ( l_23 [29] &  i[1801]);
assign l_22[24]    = ( l_23 [30] & !i[1801]) | ( l_23 [31] &  i[1801]);
assign l_22[25]    = ( l_23 [32] & !i[1801]) | ( l_23 [33] &  i[1801]);
assign l_22[26]    = ( l_23 [34]);
assign l_22[27]    = ( l_23 [35]);
assign l_23[0]    = ( l_24 [0]);
assign l_23[1]    = ( l_24 [1] & !i[1805]);
assign l_23[2]    = ( l_24 [2] & !i[1805]);
assign l_23[3]    = (!i[1805]) | ( l_24 [3] &  i[1805]);
assign l_23[4]    = (!i[1805]) | ( l_24 [4] &  i[1805]);
assign l_23[5]    = ( l_24 [5] & !i[1805]);
assign l_23[6]    = ( l_24 [6] & !i[1805]);
assign l_23[7]    = (!i[1805]) | ( l_24 [7] &  i[1805]);
assign l_23[8]    = (!i[1805]) | ( l_24 [8] &  i[1805]);
assign l_23[9]    = ( l_24 [9] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[10]    = ( l_24 [10]);
assign l_23[11]    = ( l_24 [11] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[12]    = ( l_24 [10] & !i[1805]) | ( l_24 [12] &  i[1805]);
assign l_23[13]    = ( l_24 [10] & !i[1805]) | ( l_24 [13] &  i[1805]);
assign l_23[14]    = ( l_24 [14] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[15]    = ( l_24 [15] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[16]    = ( l_24 [10] & !i[1805]) | ( l_24 [16] &  i[1805]);
assign l_23[17]    = ( l_24 [10] & !i[1805]) | ( l_24 [17] &  i[1805]);
assign l_23[18]    = ( l_24 [18] & !i[1805]) | ( l_24 [19] &  i[1805]);
assign l_23[19]    = ( l_24 [20] & !i[1805]) | ( l_24 [21] &  i[1805]);
assign l_23[20]    = ( l_24 [22] & !i[1805]) | ( l_24 [23] &  i[1805]);
assign l_23[21]    = ( l_24 [24] & !i[1805]) | ( l_24 [25] &  i[1805]);
assign l_23[22]    = ( l_24 [26] & !i[1805]) | ( l_24 [27] &  i[1805]);
assign l_23[23]    = ( l_24 [28] & !i[1805]) | ( l_24 [29] &  i[1805]);
assign l_23[24]    = ( l_24 [30] & !i[1805]) | ( l_24 [31] &  i[1805]);
assign l_23[25]    = ( l_24 [32] & !i[1805]) | ( l_24 [33] &  i[1805]);
assign l_23[26]    = ( l_24 [34] & !i[1805]) | ( l_24 [35] &  i[1805]);
assign l_23[27]    = ( l_24 [36] & !i[1805]) | ( l_24 [37] &  i[1805]);
assign l_23[28]    = ( l_24 [38] & !i[1805]) | ( l_24 [39] &  i[1805]);
assign l_23[29]    = ( l_24 [40] & !i[1805]) | ( l_24 [41] &  i[1805]);
assign l_23[30]    = ( l_24 [42] & !i[1805]) | ( l_24 [43] &  i[1805]);
assign l_23[31]    = ( l_24 [44] & !i[1805]) | ( l_24 [45] &  i[1805]);
assign l_23[32]    = ( l_24 [46] & !i[1805]) | ( l_24 [47] &  i[1805]);
assign l_23[33]    = ( l_24 [48] & !i[1805]) | ( l_24 [49] &  i[1805]);
assign l_23[34]    = ( l_24 [50]);
assign l_23[35]    = ( l_24 [51]);
assign l_24[0]    = ( l_25 [0]);
assign l_24[1]    = ( l_25 [1] & !i[1808]);
assign l_24[2]    = ( l_25 [2] & !i[1808]);
assign l_24[3]    = (!i[1808]) | ( l_25 [3] &  i[1808]);
assign l_24[4]    = (!i[1808]) | ( l_25 [4] &  i[1808]);
assign l_24[5]    = ( l_25 [5] & !i[1808]);
assign l_24[6]    = ( l_25 [6] & !i[1808]);
assign l_24[7]    = (!i[1808]) | ( l_25 [7] &  i[1808]);
assign l_24[8]    = (!i[1808]) | ( l_25 [8] &  i[1808]);
assign l_24[9]    = ( l_25 [9] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[10]    = ( l_25 [10]);
assign l_24[11]    = ( l_25 [11] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[12]    = ( l_25 [10] & !i[1808]) | ( l_25 [12] &  i[1808]);
assign l_24[13]    = ( l_25 [10] & !i[1808]) | ( l_25 [13] &  i[1808]);
assign l_24[14]    = ( l_25 [14] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[15]    = ( l_25 [15] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[16]    = ( l_25 [10] & !i[1808]) | ( l_25 [16] &  i[1808]);
assign l_24[17]    = ( l_25 [10] & !i[1808]) | ( l_25 [17] &  i[1808]);
assign l_24[18]    = ( l_25 [18]);
assign l_24[19]    = ( l_25 [19]);
assign l_24[20]    = ( l_25 [20]);
assign l_24[21]    = ( l_25 [21]);
assign l_24[22]    = ( l_25 [22]);
assign l_24[23]    = ( l_25 [23]);
assign l_24[24]    = ( l_25 [24]);
assign l_24[25]    = ( l_25 [25]);
assign l_24[26]    = ( l_25 [26]);
assign l_24[27]    = ( l_25 [27]);
assign l_24[28]    = ( l_25 [28]);
assign l_24[29]    = ( l_25 [29]);
assign l_24[30]    = ( l_25 [30]);
assign l_24[31]    = ( l_25 [31]);
assign l_24[32]    = ( l_25 [32]);
assign l_24[33]    = ( l_25 [33]);
assign l_24[34]    = ( l_25 [34]);
assign l_24[35]    = ( l_25 [35]);
assign l_24[36]    = ( l_25 [36]);
assign l_24[37]    = ( l_25 [37]);
assign l_24[38]    = ( l_25 [38]);
assign l_24[39]    = ( l_25 [39]);
assign l_24[40]    = ( l_25 [40]);
assign l_24[41]    = ( l_25 [41]);
assign l_24[42]    = ( l_25 [42]);
assign l_24[43]    = ( l_25 [43]);
assign l_24[44]    = ( l_25 [44]);
assign l_24[45]    = ( l_25 [45]);
assign l_24[46]    = ( l_25 [46]);
assign l_24[47]    = ( l_25 [47]);
assign l_24[48]    = ( l_25 [48]);
assign l_24[49]    = ( l_25 [49]);
assign l_24[50]    = ( l_25 [50] & !i[1808]) | ( l_25 [51] &  i[1808]);
assign l_24[51]    = ( l_25 [52] & !i[1808]) | ( l_25 [53] &  i[1808]);
assign l_25[0]    = ( l_26 [0]);
assign l_25[1]    = ( l_26 [1] & !i[1799]);
assign l_25[2]    = ( l_26 [2] & !i[1799]);
assign l_25[3]    = (!i[1799]) | ( l_26 [3] &  i[1799]);
assign l_25[4]    = (!i[1799]) | ( l_26 [4] &  i[1799]);
assign l_25[5]    = ( l_26 [5] & !i[1799]);
assign l_25[6]    = ( l_26 [6] & !i[1799]);
assign l_25[7]    = (!i[1799]) | ( l_26 [7] &  i[1799]);
assign l_25[8]    = (!i[1799]) | ( l_26 [8] &  i[1799]);
assign l_25[9]    = ( l_26 [9] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[10]    = ( l_26 [10]);
assign l_25[11]    = ( l_26 [11] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[12]    = ( l_26 [10] & !i[1799]) | ( l_26 [12] &  i[1799]);
assign l_25[13]    = ( l_26 [10] & !i[1799]) | ( l_26 [13] &  i[1799]);
assign l_25[14]    = ( l_26 [14] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[15]    = ( l_26 [15] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[16]    = ( l_26 [10] & !i[1799]) | ( l_26 [16] &  i[1799]);
assign l_25[17]    = ( l_26 [10] & !i[1799]) | ( l_26 [17] &  i[1799]);
assign l_25[18]    = ( l_26 [18] & !i[1799]) | ( l_26 [19] &  i[1799]);
assign l_25[19]    = ( l_26 [20] & !i[1799]) | ( l_26 [21] &  i[1799]);
assign l_25[20]    = ( l_26 [22] & !i[1799]) | ( l_26 [23] &  i[1799]);
assign l_25[21]    = ( l_26 [24] & !i[1799]) | ( l_26 [25] &  i[1799]);
assign l_25[22]    = ( l_26 [26] & !i[1799]) | ( l_26 [27] &  i[1799]);
assign l_25[23]    = ( l_26 [28] & !i[1799]) | ( l_26 [29] &  i[1799]);
assign l_25[24]    = ( l_26 [30] & !i[1799]) | ( l_26 [31] &  i[1799]);
assign l_25[25]    = ( l_26 [32] & !i[1799]) | ( l_26 [33] &  i[1799]);
assign l_25[26]    = ( l_26 [34] & !i[1799]) | ( l_26 [35] &  i[1799]);
assign l_25[27]    = ( l_26 [36] & !i[1799]) | ( l_26 [37] &  i[1799]);
assign l_25[28]    = ( l_26 [38] & !i[1799]) | ( l_26 [39] &  i[1799]);
assign l_25[29]    = ( l_26 [40] & !i[1799]) | ( l_26 [41] &  i[1799]);
assign l_25[30]    = ( l_26 [42] & !i[1799]) | ( l_26 [43] &  i[1799]);
assign l_25[31]    = ( l_26 [44] & !i[1799]) | ( l_26 [45] &  i[1799]);
assign l_25[32]    = ( l_26 [46] & !i[1799]) | ( l_26 [47] &  i[1799]);
assign l_25[33]    = ( l_26 [48] & !i[1799]) | ( l_26 [49] &  i[1799]);
assign l_25[34]    = ( l_26 [50] & !i[1799]) | ( l_26 [51] &  i[1799]);
assign l_25[35]    = ( l_26 [52] & !i[1799]) | ( l_26 [53] &  i[1799]);
assign l_25[36]    = ( l_26 [54] & !i[1799]) | ( l_26 [55] &  i[1799]);
assign l_25[37]    = ( l_26 [56] & !i[1799]) | ( l_26 [57] &  i[1799]);
assign l_25[38]    = ( l_26 [58] & !i[1799]) | ( l_26 [59] &  i[1799]);
assign l_25[39]    = ( l_26 [60] & !i[1799]) | ( l_26 [61] &  i[1799]);
assign l_25[40]    = ( l_26 [62] & !i[1799]) | ( l_26 [63] &  i[1799]);
assign l_25[41]    = ( l_26 [64] & !i[1799]) | ( l_26 [65] &  i[1799]);
assign l_25[42]    = ( l_26 [66] & !i[1799]) | ( l_26 [67] &  i[1799]);
assign l_25[43]    = ( l_26 [68] & !i[1799]) | ( l_26 [69] &  i[1799]);
assign l_25[44]    = ( l_26 [70] & !i[1799]) | ( l_26 [71] &  i[1799]);
assign l_25[45]    = ( l_26 [72] & !i[1799]) | ( l_26 [73] &  i[1799]);
assign l_25[46]    = ( l_26 [74] & !i[1799]) | ( l_26 [75] &  i[1799]);
assign l_25[47]    = ( l_26 [76] & !i[1799]) | ( l_26 [77] &  i[1799]);
assign l_25[48]    = ( l_26 [78] & !i[1799]) | ( l_26 [79] &  i[1799]);
assign l_25[49]    = ( l_26 [80] & !i[1799]) | ( l_26 [81] &  i[1799]);
assign l_25[50]    = ( l_26 [82]);
assign l_25[51]    = ( l_26 [83]);
assign l_25[52]    = ( l_26 [84]);
assign l_25[53]    = ( l_26 [85]);
assign l_26[0]    = ( l_27 [0]);
assign l_26[1]    = ( l_27 [1] & !i[1802]);
assign l_26[2]    = ( l_27 [2] & !i[1802]);
assign l_26[3]    = (!i[1802]) | ( l_27 [3] &  i[1802]);
assign l_26[4]    = (!i[1802]) | ( l_27 [4] &  i[1802]);
assign l_26[5]    = ( l_27 [5] & !i[1802]);
assign l_26[6]    = ( l_27 [6] & !i[1802]);
assign l_26[7]    = (!i[1802]) | ( l_27 [7] &  i[1802]);
assign l_26[8]    = (!i[1802]) | ( l_27 [8] &  i[1802]);
assign l_26[9]    = ( l_27 [9] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[10]    = ( l_27 [10]);
assign l_26[11]    = ( l_27 [11] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[12]    = ( l_27 [10] & !i[1802]) | ( l_27 [12] &  i[1802]);
assign l_26[13]    = ( l_27 [10] & !i[1802]) | ( l_27 [13] &  i[1802]);
assign l_26[14]    = ( l_27 [14] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[15]    = ( l_27 [15] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[16]    = ( l_27 [10] & !i[1802]) | ( l_27 [16] &  i[1802]);
assign l_26[17]    = ( l_27 [10] & !i[1802]) | ( l_27 [17] &  i[1802]);
assign l_26[18]    = ( l_27 [18]);
assign l_26[19]    = ( l_27 [19]);
assign l_26[20]    = ( l_27 [20]);
assign l_26[21]    = ( l_27 [21]);
assign l_26[22]    = ( l_27 [22]);
assign l_26[23]    = ( l_27 [23]);
assign l_26[24]    = ( l_27 [24]);
assign l_26[25]    = ( l_27 [25]);
assign l_26[26]    = ( l_27 [26]);
assign l_26[27]    = ( l_27 [27]);
assign l_26[28]    = ( l_27 [28]);
assign l_26[29]    = ( l_27 [29]);
assign l_26[30]    = ( l_27 [30]);
assign l_26[31]    = ( l_27 [31]);
assign l_26[32]    = ( l_27 [32]);
assign l_26[33]    = ( l_27 [33]);
assign l_26[34]    = ( l_27 [34]);
assign l_26[35]    = ( l_27 [35]);
assign l_26[36]    = ( l_27 [36]);
assign l_26[37]    = ( l_27 [37]);
assign l_26[38]    = ( l_27 [38]);
assign l_26[39]    = ( l_27 [39]);
assign l_26[40]    = ( l_27 [40]);
assign l_26[41]    = ( l_27 [41]);
assign l_26[42]    = ( l_27 [42]);
assign l_26[43]    = ( l_27 [43]);
assign l_26[44]    = ( l_27 [44]);
assign l_26[45]    = ( l_27 [45]);
assign l_26[46]    = ( l_27 [46]);
assign l_26[47]    = ( l_27 [47]);
assign l_26[48]    = ( l_27 [48]);
assign l_26[49]    = ( l_27 [49]);
assign l_26[50]    = ( l_27 [50]);
assign l_26[51]    = ( l_27 [51]);
assign l_26[52]    = ( l_27 [52]);
assign l_26[53]    = ( l_27 [53]);
assign l_26[54]    = ( l_27 [54]);
assign l_26[55]    = ( l_27 [55]);
assign l_26[56]    = ( l_27 [56]);
assign l_26[57]    = ( l_27 [57]);
assign l_26[58]    = ( l_27 [58]);
assign l_26[59]    = ( l_27 [59]);
assign l_26[60]    = ( l_27 [60]);
assign l_26[61]    = ( l_27 [61]);
assign l_26[62]    = ( l_27 [62]);
assign l_26[63]    = ( l_27 [63]);
assign l_26[64]    = ( l_27 [64]);
assign l_26[65]    = ( l_27 [65]);
assign l_26[66]    = ( l_27 [66]);
assign l_26[67]    = ( l_27 [67]);
assign l_26[68]    = ( l_27 [68]);
assign l_26[69]    = ( l_27 [69]);
assign l_26[70]    = ( l_27 [70]);
assign l_26[71]    = ( l_27 [71]);
assign l_26[72]    = ( l_27 [72]);
assign l_26[73]    = ( l_27 [73]);
assign l_26[74]    = ( l_27 [74]);
assign l_26[75]    = ( l_27 [75]);
assign l_26[76]    = ( l_27 [76]);
assign l_26[77]    = ( l_27 [77]);
assign l_26[78]    = ( l_27 [78]);
assign l_26[79]    = ( l_27 [79]);
assign l_26[80]    = ( l_27 [80]);
assign l_26[81]    = ( l_27 [81]);
assign l_26[82]    = ( l_27 [82] & !i[1802]) | ( l_27 [83] &  i[1802]);
assign l_26[83]    = ( l_27 [84] & !i[1802]) | ( l_27 [85] &  i[1802]);
assign l_26[84]    = ( l_27 [86] & !i[1802]) | ( l_27 [87] &  i[1802]);
assign l_26[85]    = ( l_27 [88] & !i[1802]) | ( l_27 [89] &  i[1802]);
assign l_27[0]    = ( l_28 [0]);
assign l_27[1]    = ( l_28 [1] & !i[1806]);
assign l_27[2]    = ( l_28 [2] & !i[1806]);
assign l_27[3]    = (!i[1806]) | ( l_28 [3] &  i[1806]);
assign l_27[4]    = (!i[1806]) | ( l_28 [4] &  i[1806]);
assign l_27[5]    = ( l_28 [5] & !i[1806]);
assign l_27[6]    = ( l_28 [6] & !i[1806]);
assign l_27[7]    = (!i[1806]) | ( l_28 [7] &  i[1806]);
assign l_27[8]    = (!i[1806]) | ( l_28 [8] &  i[1806]);
assign l_27[9]    = ( l_28 [9] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[10]    = ( l_28 [10]);
assign l_27[11]    = ( l_28 [11] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[12]    = ( l_28 [10] & !i[1806]) | ( l_28 [12] &  i[1806]);
assign l_27[13]    = ( l_28 [10] & !i[1806]) | ( l_28 [13] &  i[1806]);
assign l_27[14]    = ( l_28 [14] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[15]    = ( l_28 [15] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[16]    = ( l_28 [10] & !i[1806]) | ( l_28 [16] &  i[1806]);
assign l_27[17]    = ( l_28 [10] & !i[1806]) | ( l_28 [17] &  i[1806]);
assign l_27[18]    = ( l_28 [18]);
assign l_27[19]    = ( l_28 [19]);
assign l_27[20]    = ( l_28 [20]);
assign l_27[21]    = ( l_28 [21]);
assign l_27[22]    = ( l_28 [22]);
assign l_27[23]    = ( l_28 [23]);
assign l_27[24]    = ( l_28 [24]);
assign l_27[25]    = ( l_28 [25]);
assign l_27[26]    = ( l_28 [26]);
assign l_27[27]    = ( l_28 [27]);
assign l_27[28]    = ( l_28 [28]);
assign l_27[29]    = ( l_28 [29]);
assign l_27[30]    = ( l_28 [30]);
assign l_27[31]    = ( l_28 [31]);
assign l_27[32]    = ( l_28 [32]);
assign l_27[33]    = ( l_28 [33]);
assign l_27[34]    = ( l_28 [34]);
assign l_27[35]    = ( l_28 [35]);
assign l_27[36]    = ( l_28 [36]);
assign l_27[37]    = ( l_28 [37]);
assign l_27[38]    = ( l_28 [38]);
assign l_27[39]    = ( l_28 [39]);
assign l_27[40]    = ( l_28 [40]);
assign l_27[41]    = ( l_28 [41]);
assign l_27[42]    = ( l_28 [42]);
assign l_27[43]    = ( l_28 [43]);
assign l_27[44]    = ( l_28 [44]);
assign l_27[45]    = ( l_28 [45]);
assign l_27[46]    = ( l_28 [46]);
assign l_27[47]    = ( l_28 [47]);
assign l_27[48]    = ( l_28 [48]);
assign l_27[49]    = ( l_28 [49]);
assign l_27[50]    = ( l_28 [50]);
assign l_27[51]    = ( l_28 [51]);
assign l_27[52]    = ( l_28 [52]);
assign l_27[53]    = ( l_28 [53]);
assign l_27[54]    = ( l_28 [54]);
assign l_27[55]    = ( l_28 [55]);
assign l_27[56]    = ( l_28 [56]);
assign l_27[57]    = ( l_28 [57]);
assign l_27[58]    = ( l_28 [58]);
assign l_27[59]    = ( l_28 [59]);
assign l_27[60]    = ( l_28 [60]);
assign l_27[61]    = ( l_28 [61]);
assign l_27[62]    = ( l_28 [62]);
assign l_27[63]    = ( l_28 [63]);
assign l_27[64]    = ( l_28 [64]);
assign l_27[65]    = ( l_28 [65]);
assign l_27[66]    = ( l_28 [66]);
assign l_27[67]    = ( l_28 [67]);
assign l_27[68]    = ( l_28 [68]);
assign l_27[69]    = ( l_28 [69]);
assign l_27[70]    = ( l_28 [70]);
assign l_27[71]    = ( l_28 [71]);
assign l_27[72]    = ( l_28 [72]);
assign l_27[73]    = ( l_28 [73]);
assign l_27[74]    = ( l_28 [74]);
assign l_27[75]    = ( l_28 [75]);
assign l_27[76]    = ( l_28 [76]);
assign l_27[77]    = ( l_28 [77]);
assign l_27[78]    = ( l_28 [78]);
assign l_27[79]    = ( l_28 [79]);
assign l_27[80]    = ( l_28 [80]);
assign l_27[81]    = ( l_28 [81]);
assign l_27[82]    = ( l_28 [82] & !i[1806]) | ( l_28 [83] &  i[1806]);
assign l_27[83]    = ( l_28 [84] & !i[1806]) | ( l_28 [85] &  i[1806]);
assign l_27[84]    = ( l_28 [86] & !i[1806]) | ( l_28 [87] &  i[1806]);
assign l_27[85]    = ( l_28 [88] & !i[1806]) | ( l_28 [89] &  i[1806]);
assign l_27[86]    = ( l_28 [90] & !i[1806]) | ( l_28 [91] &  i[1806]);
assign l_27[87]    = ( l_28 [92] & !i[1806]) | ( l_28 [93] &  i[1806]);
assign l_27[88]    = ( l_28 [94] & !i[1806]) | ( l_28 [95] &  i[1806]);
assign l_27[89]    = ( l_28 [96] & !i[1806]) | ( l_28 [97] &  i[1806]);
assign l_28[0]    = ( l_29 [0]);
assign l_28[1]    = ( l_29 [1] & !i[1816]);
assign l_28[2]    = ( l_29 [2] & !i[1816]);
assign l_28[3]    = (!i[1816]) | ( l_29 [3] &  i[1816]);
assign l_28[4]    = (!i[1816]) | ( l_29 [4] &  i[1816]);
assign l_28[5]    = ( l_29 [5] & !i[1816]);
assign l_28[6]    = ( l_29 [6] & !i[1816]);
assign l_28[7]    = (!i[1816]) | ( l_29 [7] &  i[1816]);
assign l_28[8]    = (!i[1816]) | ( l_29 [8] &  i[1816]);
assign l_28[9]    = ( l_29 [9] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[10]    = ( l_29 [10]);
assign l_28[11]    = ( l_29 [11] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[12]    = ( l_29 [10] & !i[1816]) | ( l_29 [12] &  i[1816]);
assign l_28[13]    = ( l_29 [10] & !i[1816]) | ( l_29 [13] &  i[1816]);
assign l_28[14]    = ( l_29 [14] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[15]    = ( l_29 [15] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[16]    = ( l_29 [10] & !i[1816]) | ( l_29 [16] &  i[1816]);
assign l_28[17]    = ( l_29 [10] & !i[1816]) | ( l_29 [17] &  i[1816]);
assign l_28[18]    = ( l_29 [18]);
assign l_28[19]    = ( l_29 [19]);
assign l_28[20]    = ( l_29 [20]);
assign l_28[21]    = ( l_29 [21]);
assign l_28[22]    = ( l_29 [22]);
assign l_28[23]    = ( l_29 [23]);
assign l_28[24]    = ( l_29 [24]);
assign l_28[25]    = ( l_29 [25]);
assign l_28[26]    = ( l_29 [26]);
assign l_28[27]    = ( l_29 [27]);
assign l_28[28]    = ( l_29 [28]);
assign l_28[29]    = ( l_29 [29]);
assign l_28[30]    = ( l_29 [30]);
assign l_28[31]    = ( l_29 [31]);
assign l_28[32]    = ( l_29 [32]);
assign l_28[33]    = ( l_29 [33]);
assign l_28[34]    = ( l_29 [34]);
assign l_28[35]    = ( l_29 [35]);
assign l_28[36]    = ( l_29 [36]);
assign l_28[37]    = ( l_29 [37]);
assign l_28[38]    = ( l_29 [38]);
assign l_28[39]    = ( l_29 [39]);
assign l_28[40]    = ( l_29 [40]);
assign l_28[41]    = ( l_29 [41]);
assign l_28[42]    = ( l_29 [42]);
assign l_28[43]    = ( l_29 [43]);
assign l_28[44]    = ( l_29 [44]);
assign l_28[45]    = ( l_29 [45]);
assign l_28[46]    = ( l_29 [46]);
assign l_28[47]    = ( l_29 [47]);
assign l_28[48]    = ( l_29 [48]);
assign l_28[49]    = ( l_29 [49]);
assign l_28[50]    = ( l_29 [50]);
assign l_28[51]    = ( l_29 [51]);
assign l_28[52]    = ( l_29 [52]);
assign l_28[53]    = ( l_29 [53]);
assign l_28[54]    = ( l_29 [54]);
assign l_28[55]    = ( l_29 [55]);
assign l_28[56]    = ( l_29 [56]);
assign l_28[57]    = ( l_29 [57]);
assign l_28[58]    = ( l_29 [58]);
assign l_28[59]    = ( l_29 [59]);
assign l_28[60]    = ( l_29 [60]);
assign l_28[61]    = ( l_29 [61]);
assign l_28[62]    = ( l_29 [62]);
assign l_28[63]    = ( l_29 [63]);
assign l_28[64]    = ( l_29 [64]);
assign l_28[65]    = ( l_29 [65]);
assign l_28[66]    = ( l_29 [66]);
assign l_28[67]    = ( l_29 [67]);
assign l_28[68]    = ( l_29 [68]);
assign l_28[69]    = ( l_29 [69]);
assign l_28[70]    = ( l_29 [70]);
assign l_28[71]    = ( l_29 [71]);
assign l_28[72]    = ( l_29 [72]);
assign l_28[73]    = ( l_29 [73]);
assign l_28[74]    = ( l_29 [74]);
assign l_28[75]    = ( l_29 [75]);
assign l_28[76]    = ( l_29 [76]);
assign l_28[77]    = ( l_29 [77]);
assign l_28[78]    = ( l_29 [78]);
assign l_28[79]    = ( l_29 [79]);
assign l_28[80]    = ( l_29 [80]);
assign l_28[81]    = ( l_29 [81]);
assign l_28[82]    = ( l_29 [82] & !i[1816]) | ( l_29 [83] &  i[1816]);
assign l_28[83]    = ( l_29 [84] & !i[1816]) | ( l_29 [85] &  i[1816]);
assign l_28[84]    = ( l_29 [86] & !i[1816]) | ( l_29 [87] &  i[1816]);
assign l_28[85]    = ( l_29 [88] & !i[1816]) | ( l_29 [89] &  i[1816]);
assign l_28[86]    = ( l_29 [90] & !i[1816]) | ( l_29 [91] &  i[1816]);
assign l_28[87]    = ( l_29 [92] & !i[1816]) | ( l_29 [93] &  i[1816]);
assign l_28[88]    = ( l_29 [94] & !i[1816]) | ( l_29 [95] &  i[1816]);
assign l_28[89]    = ( l_29 [96] & !i[1816]) | ( l_29 [97] &  i[1816]);
assign l_28[90]    = ( l_29 [98] & !i[1816]) | ( l_29 [99] &  i[1816]);
assign l_28[91]    = ( l_29 [100] & !i[1816]) | ( l_29 [101] &  i[1816]);
assign l_28[92]    = ( l_29 [102] & !i[1816]) | ( l_29 [103] &  i[1816]);
assign l_28[93]    = ( l_29 [104] & !i[1816]) | ( l_29 [105] &  i[1816]);
assign l_28[94]    = ( l_29 [106] & !i[1816]) | ( l_29 [107] &  i[1816]);
assign l_28[95]    = ( l_29 [108] & !i[1816]) | ( l_29 [109] &  i[1816]);
assign l_28[96]    = ( l_29 [110] & !i[1816]) | ( l_29 [111] &  i[1816]);
assign l_28[97]    = ( l_29 [112] & !i[1816]) | ( l_29 [113] &  i[1816]);
assign l_29[0]    = ( l_30 [0]);
assign l_29[1]    = ( l_30 [1] & !i[1810]);
assign l_29[2]    = ( l_30 [2] & !i[1810]);
assign l_29[3]    = (!i[1810]) | ( l_30 [3] &  i[1810]);
assign l_29[4]    = (!i[1810]) | ( l_30 [4] &  i[1810]);
assign l_29[5]    = ( l_30 [5] & !i[1810]);
assign l_29[6]    = ( l_30 [6] & !i[1810]);
assign l_29[7]    = (!i[1810]) | ( l_30 [7] &  i[1810]);
assign l_29[8]    = (!i[1810]) | ( l_30 [8] &  i[1810]);
assign l_29[9]    = ( l_30 [9] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[10]    = ( l_30 [10]);
assign l_29[11]    = ( l_30 [11] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[12]    = ( l_30 [10] & !i[1810]) | ( l_30 [12] &  i[1810]);
assign l_29[13]    = ( l_30 [10] & !i[1810]) | ( l_30 [13] &  i[1810]);
assign l_29[14]    = ( l_30 [14] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[15]    = ( l_30 [15] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[16]    = ( l_30 [10] & !i[1810]) | ( l_30 [16] &  i[1810]);
assign l_29[17]    = ( l_30 [10] & !i[1810]) | ( l_30 [17] &  i[1810]);
assign l_29[18]    = ( l_30 [18]);
assign l_29[19]    = ( l_30 [19]);
assign l_29[20]    = ( l_30 [20]);
assign l_29[21]    = ( l_30 [21]);
assign l_29[22]    = ( l_30 [22]);
assign l_29[23]    = ( l_30 [23]);
assign l_29[24]    = ( l_30 [24]);
assign l_29[25]    = ( l_30 [25]);
assign l_29[26]    = ( l_30 [26]);
assign l_29[27]    = ( l_30 [27]);
assign l_29[28]    = ( l_30 [28]);
assign l_29[29]    = ( l_30 [29]);
assign l_29[30]    = ( l_30 [30]);
assign l_29[31]    = ( l_30 [31]);
assign l_29[32]    = ( l_30 [32]);
assign l_29[33]    = ( l_30 [33]);
assign l_29[34]    = ( l_30 [34]);
assign l_29[35]    = ( l_30 [35]);
assign l_29[36]    = ( l_30 [36]);
assign l_29[37]    = ( l_30 [37]);
assign l_29[38]    = ( l_30 [38]);
assign l_29[39]    = ( l_30 [39]);
assign l_29[40]    = ( l_30 [40]);
assign l_29[41]    = ( l_30 [41]);
assign l_29[42]    = ( l_30 [42]);
assign l_29[43]    = ( l_30 [43]);
assign l_29[44]    = ( l_30 [44]);
assign l_29[45]    = ( l_30 [45]);
assign l_29[46]    = ( l_30 [46]);
assign l_29[47]    = ( l_30 [47]);
assign l_29[48]    = ( l_30 [48]);
assign l_29[49]    = ( l_30 [49]);
assign l_29[50]    = ( l_30 [50]);
assign l_29[51]    = ( l_30 [51]);
assign l_29[52]    = ( l_30 [52]);
assign l_29[53]    = ( l_30 [53]);
assign l_29[54]    = ( l_30 [54]);
assign l_29[55]    = ( l_30 [55]);
assign l_29[56]    = ( l_30 [56]);
assign l_29[57]    = ( l_30 [57]);
assign l_29[58]    = ( l_30 [58]);
assign l_29[59]    = ( l_30 [59]);
assign l_29[60]    = ( l_30 [60]);
assign l_29[61]    = ( l_30 [61]);
assign l_29[62]    = ( l_30 [62]);
assign l_29[63]    = ( l_30 [63]);
assign l_29[64]    = ( l_30 [64]);
assign l_29[65]    = ( l_30 [65]);
assign l_29[66]    = ( l_30 [66]);
assign l_29[67]    = ( l_30 [67]);
assign l_29[68]    = ( l_30 [68]);
assign l_29[69]    = ( l_30 [69]);
assign l_29[70]    = ( l_30 [70]);
assign l_29[71]    = ( l_30 [71]);
assign l_29[72]    = ( l_30 [72]);
assign l_29[73]    = ( l_30 [73]);
assign l_29[74]    = ( l_30 [74]);
assign l_29[75]    = ( l_30 [75]);
assign l_29[76]    = ( l_30 [76]);
assign l_29[77]    = ( l_30 [77]);
assign l_29[78]    = ( l_30 [78]);
assign l_29[79]    = ( l_30 [79]);
assign l_29[80]    = ( l_30 [80]);
assign l_29[81]    = ( l_30 [81]);
assign l_29[82]    = ( l_30 [82] & !i[1810]) | ( l_30 [83] &  i[1810]);
assign l_29[83]    = ( l_30 [84] & !i[1810]) | ( l_30 [85] &  i[1810]);
assign l_29[84]    = ( l_30 [86] & !i[1810]) | ( l_30 [87] &  i[1810]);
assign l_29[85]    = ( l_30 [88] & !i[1810]) | ( l_30 [89] &  i[1810]);
assign l_29[86]    = ( l_30 [90] & !i[1810]) | ( l_30 [91] &  i[1810]);
assign l_29[87]    = ( l_30 [92] & !i[1810]) | ( l_30 [93] &  i[1810]);
assign l_29[88]    = ( l_30 [94] & !i[1810]) | ( l_30 [95] &  i[1810]);
assign l_29[89]    = ( l_30 [96] & !i[1810]) | ( l_30 [97] &  i[1810]);
assign l_29[90]    = ( l_30 [98] & !i[1810]) | ( l_30 [99] &  i[1810]);
assign l_29[91]    = ( l_30 [100] & !i[1810]) | ( l_30 [101] &  i[1810]);
assign l_29[92]    = ( l_30 [102] & !i[1810]) | ( l_30 [103] &  i[1810]);
assign l_29[93]    = ( l_30 [104] & !i[1810]) | ( l_30 [105] &  i[1810]);
assign l_29[94]    = ( l_30 [106] & !i[1810]) | ( l_30 [107] &  i[1810]);
assign l_29[95]    = ( l_30 [108] & !i[1810]) | ( l_30 [109] &  i[1810]);
assign l_29[96]    = ( l_30 [110] & !i[1810]) | ( l_30 [111] &  i[1810]);
assign l_29[97]    = ( l_30 [112] & !i[1810]) | ( l_30 [113] &  i[1810]);
assign l_29[98]    = ( l_30 [114] & !i[1810]) | ( l_30 [115] &  i[1810]);
assign l_29[99]    = ( l_30 [116] & !i[1810]) | ( l_30 [117] &  i[1810]);
assign l_29[100]    = ( l_30 [118] & !i[1810]) | ( l_30 [119] &  i[1810]);
assign l_29[101]    = ( l_30 [120] & !i[1810]) | ( l_30 [121] &  i[1810]);
assign l_29[102]    = ( l_30 [122] & !i[1810]) | ( l_30 [123] &  i[1810]);
assign l_29[103]    = ( l_30 [124] & !i[1810]) | ( l_30 [125] &  i[1810]);
assign l_29[104]    = ( l_30 [126] & !i[1810]) | ( l_30 [127] &  i[1810]);
assign l_29[105]    = ( l_30 [128] & !i[1810]) | ( l_30 [129] &  i[1810]);
assign l_29[106]    = ( l_30 [130] & !i[1810]) | ( l_30 [131] &  i[1810]);
assign l_29[107]    = ( l_30 [132] & !i[1810]) | ( l_30 [133] &  i[1810]);
assign l_29[108]    = ( l_30 [134] & !i[1810]) | ( l_30 [135] &  i[1810]);
assign l_29[109]    = ( l_30 [136] & !i[1810]) | ( l_30 [137] &  i[1810]);
assign l_29[110]    = ( l_30 [138] & !i[1810]) | ( l_30 [139] &  i[1810]);
assign l_29[111]    = ( l_30 [140] & !i[1810]) | ( l_30 [141] &  i[1810]);
assign l_29[112]    = ( l_30 [142] & !i[1810]) | ( l_30 [143] &  i[1810]);
assign l_29[113]    = ( l_30 [144] & !i[1810]) | ( l_30 [145] &  i[1810]);
assign l_30[0]    = ( l_31 [0]);
assign l_30[1]    = ( l_31 [1] & !i[1804]);
assign l_30[2]    = ( l_31 [2] & !i[1804]);
assign l_30[3]    = (!i[1804]) | ( l_31 [3] &  i[1804]);
assign l_30[4]    = (!i[1804]) | ( l_31 [4] &  i[1804]);
assign l_30[5]    = ( l_31 [5] & !i[1804]);
assign l_30[6]    = ( l_31 [6] & !i[1804]);
assign l_30[7]    = (!i[1804]) | ( l_31 [7] &  i[1804]);
assign l_30[8]    = (!i[1804]) | ( l_31 [8] &  i[1804]);
assign l_30[9]    = ( l_31 [9] & !i[1804]) | ( l_31 [10] &  i[1804]);
assign l_30[10]    = ( l_31 [10]);
assign l_30[11]    = ( l_31 [11] & !i[1804]) | ( l_31 [10] &  i[1804]);
assign l_30[12]    = ( l_31 [10] & !i[1804]) | ( l_31 [12] &  i[1804]);
assign l_30[13]    = ( l_31 [10] & !i[1804]) | ( l_31 [13] &  i[1804]);
assign l_30[14]    = ( l_31 [14] & !i[1804]) | ( l_31 [10] &  i[1804]);
assign l_30[15]    = ( l_31 [15] & !i[1804]) | ( l_31 [10] &  i[1804]);
assign l_30[16]    = ( l_31 [10] & !i[1804]) | ( l_31 [16] &  i[1804]);
assign l_30[17]    = ( l_31 [10] & !i[1804]) | ( l_31 [17] &  i[1804]);
assign l_30[18]    = ( l_31 [18]);
assign l_30[19]    = ( l_31 [19]);
assign l_30[20]    = ( l_31 [20]);
assign l_30[21]    = ( l_31 [21]);
assign l_30[22]    = ( l_31 [22]);
assign l_30[23]    = ( l_31 [23]);
assign l_30[24]    = ( l_31 [24]);
assign l_30[25]    = ( l_31 [25]);
assign l_30[26]    = ( l_31 [26]);
assign l_30[27]    = ( l_31 [27]);
assign l_30[28]    = ( l_31 [28]);
assign l_30[29]    = ( l_31 [29]);
assign l_30[30]    = ( l_31 [30]);
assign l_30[31]    = ( l_31 [31]);
assign l_30[32]    = ( l_31 [32]);
assign l_30[33]    = ( l_31 [33]);
assign l_30[34]    = ( l_31 [34]);
assign l_30[35]    = ( l_31 [35]);
assign l_30[36]    = ( l_31 [36]);
assign l_30[37]    = ( l_31 [37]);
assign l_30[38]    = ( l_31 [38]);
assign l_30[39]    = ( l_31 [39]);
assign l_30[40]    = ( l_31 [40]);
assign l_30[41]    = ( l_31 [41]);
assign l_30[42]    = ( l_31 [42]);
assign l_30[43]    = ( l_31 [43]);
assign l_30[44]    = ( l_31 [44]);
assign l_30[45]    = ( l_31 [45]);
assign l_30[46]    = ( l_31 [46]);
assign l_30[47]    = ( l_31 [47]);
assign l_30[48]    = ( l_31 [48]);
assign l_30[49]    = ( l_31 [49]);
assign l_30[50]    = ( l_31 [50]);
assign l_30[51]    = ( l_31 [51]);
assign l_30[52]    = ( l_31 [52]);
assign l_30[53]    = ( l_31 [53]);
assign l_30[54]    = ( l_31 [54]);
assign l_30[55]    = ( l_31 [55]);
assign l_30[56]    = ( l_31 [56]);
assign l_30[57]    = ( l_31 [57]);
assign l_30[58]    = ( l_31 [58]);
assign l_30[59]    = ( l_31 [59]);
assign l_30[60]    = ( l_31 [60]);
assign l_30[61]    = ( l_31 [61]);
assign l_30[62]    = ( l_31 [62]);
assign l_30[63]    = ( l_31 [63]);
assign l_30[64]    = ( l_31 [64]);
assign l_30[65]    = ( l_31 [65]);
assign l_30[66]    = ( l_31 [66]);
assign l_30[67]    = ( l_31 [67]);
assign l_30[68]    = ( l_31 [68]);
assign l_30[69]    = ( l_31 [69]);
assign l_30[70]    = ( l_31 [70]);
assign l_30[71]    = ( l_31 [71]);
assign l_30[72]    = ( l_31 [72]);
assign l_30[73]    = ( l_31 [73]);
assign l_30[74]    = ( l_31 [74]);
assign l_30[75]    = ( l_31 [75]);
assign l_30[76]    = ( l_31 [76]);
assign l_30[77]    = ( l_31 [77]);
assign l_30[78]    = ( l_31 [78]);
assign l_30[79]    = ( l_31 [79]);
assign l_30[80]    = ( l_31 [80]);
assign l_30[81]    = ( l_31 [81]);
assign l_30[82]    = ( l_31 [82] & !i[1804]) | ( l_31 [83] &  i[1804]);
assign l_30[83]    = ( l_31 [84] & !i[1804]) | ( l_31 [85] &  i[1804]);
assign l_30[84]    = ( l_31 [86] & !i[1804]) | ( l_31 [87] &  i[1804]);
assign l_30[85]    = ( l_31 [88] & !i[1804]) | ( l_31 [89] &  i[1804]);
assign l_30[86]    = ( l_31 [90] & !i[1804]) | ( l_31 [91] &  i[1804]);
assign l_30[87]    = ( l_31 [92] & !i[1804]) | ( l_31 [93] &  i[1804]);
assign l_30[88]    = ( l_31 [94] & !i[1804]) | ( l_31 [95] &  i[1804]);
assign l_30[89]    = ( l_31 [96] & !i[1804]) | ( l_31 [97] &  i[1804]);
assign l_30[90]    = ( l_31 [98] & !i[1804]) | ( l_31 [99] &  i[1804]);
assign l_30[91]    = ( l_31 [100] & !i[1804]) | ( l_31 [101] &  i[1804]);
assign l_30[92]    = ( l_31 [102] & !i[1804]) | ( l_31 [103] &  i[1804]);
assign l_30[93]    = ( l_31 [104] & !i[1804]) | ( l_31 [105] &  i[1804]);
assign l_30[94]    = ( l_31 [106] & !i[1804]) | ( l_31 [107] &  i[1804]);
assign l_30[95]    = ( l_31 [108] & !i[1804]) | ( l_31 [109] &  i[1804]);
assign l_30[96]    = ( l_31 [110] & !i[1804]) | ( l_31 [111] &  i[1804]);
assign l_30[97]    = ( l_31 [112] & !i[1804]) | ( l_31 [113] &  i[1804]);
assign l_30[98]    = ( l_31 [114] & !i[1804]) | ( l_31 [115] &  i[1804]);
assign l_30[99]    = ( l_31 [116] & !i[1804]) | ( l_31 [117] &  i[1804]);
assign l_30[100]    = ( l_31 [118] & !i[1804]) | ( l_31 [119] &  i[1804]);
assign l_30[101]    = ( l_31 [120] & !i[1804]) | ( l_31 [121] &  i[1804]);
assign l_30[102]    = ( l_31 [122] & !i[1804]) | ( l_31 [123] &  i[1804]);
assign l_30[103]    = ( l_31 [124] & !i[1804]) | ( l_31 [125] &  i[1804]);
assign l_30[104]    = ( l_31 [126] & !i[1804]) | ( l_31 [127] &  i[1804]);
assign l_30[105]    = ( l_31 [128] & !i[1804]) | ( l_31 [129] &  i[1804]);
assign l_30[106]    = ( l_31 [130] & !i[1804]) | ( l_31 [131] &  i[1804]);
assign l_30[107]    = ( l_31 [132] & !i[1804]) | ( l_31 [133] &  i[1804]);
assign l_30[108]    = ( l_31 [134] & !i[1804]) | ( l_31 [135] &  i[1804]);
assign l_30[109]    = ( l_31 [136] & !i[1804]) | ( l_31 [137] &  i[1804]);
assign l_30[110]    = ( l_31 [138] & !i[1804]) | ( l_31 [139] &  i[1804]);
assign l_30[111]    = ( l_31 [140] & !i[1804]) | ( l_31 [141] &  i[1804]);
assign l_30[112]    = ( l_31 [142] & !i[1804]) | ( l_31 [143] &  i[1804]);
assign l_30[113]    = ( l_31 [144] & !i[1804]) | ( l_31 [145] &  i[1804]);
assign l_30[114]    = ( l_31 [146] & !i[1804]) | ( l_31 [147] &  i[1804]);
assign l_30[115]    = ( l_31 [148] & !i[1804]) | ( l_31 [149] &  i[1804]);
assign l_30[116]    = ( l_31 [150] & !i[1804]) | ( l_31 [151] &  i[1804]);
assign l_30[117]    = ( l_31 [152] & !i[1804]) | ( l_31 [153] &  i[1804]);
assign l_30[118]    = ( l_31 [154] & !i[1804]) | ( l_31 [155] &  i[1804]);
assign l_30[119]    = ( l_31 [156] & !i[1804]) | ( l_31 [157] &  i[1804]);
assign l_30[120]    = ( l_31 [158] & !i[1804]) | ( l_31 [159] &  i[1804]);
assign l_30[121]    = ( l_31 [160] & !i[1804]) | ( l_31 [161] &  i[1804]);
assign l_30[122]    = ( l_31 [162] & !i[1804]) | ( l_31 [163] &  i[1804]);
assign l_30[123]    = ( l_31 [164] & !i[1804]) | ( l_31 [165] &  i[1804]);
assign l_30[124]    = ( l_31 [166] & !i[1804]) | ( l_31 [167] &  i[1804]);
assign l_30[125]    = ( l_31 [168] & !i[1804]) | ( l_31 [169] &  i[1804]);
assign l_30[126]    = ( l_31 [170] & !i[1804]) | ( l_31 [171] &  i[1804]);
assign l_30[127]    = ( l_31 [172] & !i[1804]) | ( l_31 [173] &  i[1804]);
assign l_30[128]    = ( l_31 [174] & !i[1804]) | ( l_31 [175] &  i[1804]);
assign l_30[129]    = ( l_31 [176] & !i[1804]) | ( l_31 [177] &  i[1804]);
assign l_30[130]    = ( l_31 [178] & !i[1804]) | ( l_31 [179] &  i[1804]);
assign l_30[131]    = ( l_31 [180] & !i[1804]) | ( l_31 [181] &  i[1804]);
assign l_30[132]    = ( l_31 [182] & !i[1804]) | ( l_31 [183] &  i[1804]);
assign l_30[133]    = ( l_31 [184] & !i[1804]) | ( l_31 [185] &  i[1804]);
assign l_30[134]    = ( l_31 [186] & !i[1804]) | ( l_31 [187] &  i[1804]);
assign l_30[135]    = ( l_31 [188] & !i[1804]) | ( l_31 [189] &  i[1804]);
assign l_30[136]    = ( l_31 [190] & !i[1804]) | ( l_31 [191] &  i[1804]);
assign l_30[137]    = ( l_31 [192] & !i[1804]) | ( l_31 [193] &  i[1804]);
assign l_30[138]    = ( l_31 [194] & !i[1804]) | ( l_31 [195] &  i[1804]);
assign l_30[139]    = ( l_31 [196] & !i[1804]) | ( l_31 [197] &  i[1804]);
assign l_30[140]    = ( l_31 [198] & !i[1804]) | ( l_31 [199] &  i[1804]);
assign l_30[141]    = ( l_31 [200] & !i[1804]) | ( l_31 [201] &  i[1804]);
assign l_30[142]    = ( l_31 [202] & !i[1804]) | ( l_31 [203] &  i[1804]);
assign l_30[143]    = ( l_31 [204] & !i[1804]) | ( l_31 [205] &  i[1804]);
assign l_30[144]    = ( l_31 [206] & !i[1804]) | ( l_31 [207] &  i[1804]);
assign l_30[145]    = ( l_31 [208] & !i[1804]) | ( l_31 [209] &  i[1804]);
assign l_31[0]    = ( l_32 [0]);
assign l_31[1]    = ( l_32 [1] & !i[1811]);
assign l_31[2]    = ( l_32 [2] & !i[1811]);
assign l_31[3]    = (!i[1811]) | ( l_32 [3] &  i[1811]);
assign l_31[4]    = (!i[1811]) | ( l_32 [4] &  i[1811]);
assign l_31[5]    = ( l_32 [5] & !i[1811]);
assign l_31[6]    = ( l_32 [6] & !i[1811]);
assign l_31[7]    = (!i[1811]) | ( l_32 [7] &  i[1811]);
assign l_31[8]    = (!i[1811]) | ( l_32 [8] &  i[1811]);
assign l_31[9]    = ( l_32 [9] & !i[1811]) | ( l_32 [10] &  i[1811]);
assign l_31[10]    = ( l_32 [10]);
assign l_31[11]    = ( l_32 [11] & !i[1811]) | ( l_32 [10] &  i[1811]);
assign l_31[12]    = ( l_32 [10] & !i[1811]) | ( l_32 [12] &  i[1811]);
assign l_31[13]    = ( l_32 [10] & !i[1811]) | ( l_32 [13] &  i[1811]);
assign l_31[14]    = ( l_32 [14] & !i[1811]) | ( l_32 [10] &  i[1811]);
assign l_31[15]    = ( l_32 [15] & !i[1811]) | ( l_32 [10] &  i[1811]);
assign l_31[16]    = ( l_32 [10] & !i[1811]) | ( l_32 [16] &  i[1811]);
assign l_31[17]    = ( l_32 [10] & !i[1811]) | ( l_32 [17] &  i[1811]);
assign l_31[18]    = ( l_32 [18] & !i[1811]) | ( l_32 [19] &  i[1811]);
assign l_31[19]    = ( l_32 [20] & !i[1811]) | ( l_32 [21] &  i[1811]);
assign l_31[20]    = ( l_32 [22] & !i[1811]) | ( l_32 [23] &  i[1811]);
assign l_31[21]    = ( l_32 [24] & !i[1811]) | ( l_32 [25] &  i[1811]);
assign l_31[22]    = ( l_32 [26] & !i[1811]) | ( l_32 [27] &  i[1811]);
assign l_31[23]    = ( l_32 [28] & !i[1811]) | ( l_32 [29] &  i[1811]);
assign l_31[24]    = ( l_32 [30] & !i[1811]) | ( l_32 [31] &  i[1811]);
assign l_31[25]    = ( l_32 [32] & !i[1811]) | ( l_32 [33] &  i[1811]);
assign l_31[26]    = ( l_32 [34] & !i[1811]) | ( l_32 [35] &  i[1811]);
assign l_31[27]    = ( l_32 [36] & !i[1811]) | ( l_32 [37] &  i[1811]);
assign l_31[28]    = ( l_32 [38] & !i[1811]) | ( l_32 [39] &  i[1811]);
assign l_31[29]    = ( l_32 [40] & !i[1811]) | ( l_32 [41] &  i[1811]);
assign l_31[30]    = ( l_32 [42] & !i[1811]) | ( l_32 [43] &  i[1811]);
assign l_31[31]    = ( l_32 [44] & !i[1811]) | ( l_32 [45] &  i[1811]);
assign l_31[32]    = ( l_32 [46] & !i[1811]) | ( l_32 [47] &  i[1811]);
assign l_31[33]    = ( l_32 [48] & !i[1811]) | ( l_32 [49] &  i[1811]);
assign l_31[34]    = ( l_32 [50] & !i[1811]) | ( l_32 [51] &  i[1811]);
assign l_31[35]    = ( l_32 [52] & !i[1811]) | ( l_32 [53] &  i[1811]);
assign l_31[36]    = ( l_32 [54] & !i[1811]) | ( l_32 [55] &  i[1811]);
assign l_31[37]    = ( l_32 [56] & !i[1811]) | ( l_32 [57] &  i[1811]);
assign l_31[38]    = ( l_32 [58] & !i[1811]) | ( l_32 [59] &  i[1811]);
assign l_31[39]    = ( l_32 [60] & !i[1811]) | ( l_32 [61] &  i[1811]);
assign l_31[40]    = ( l_32 [62] & !i[1811]) | ( l_32 [63] &  i[1811]);
assign l_31[41]    = ( l_32 [64] & !i[1811]) | ( l_32 [65] &  i[1811]);
assign l_31[42]    = ( l_32 [66] & !i[1811]) | ( l_32 [67] &  i[1811]);
assign l_31[43]    = ( l_32 [68] & !i[1811]) | ( l_32 [69] &  i[1811]);
assign l_31[44]    = ( l_32 [70] & !i[1811]) | ( l_32 [71] &  i[1811]);
assign l_31[45]    = ( l_32 [72] & !i[1811]) | ( l_32 [73] &  i[1811]);
assign l_31[46]    = ( l_32 [74] & !i[1811]) | ( l_32 [75] &  i[1811]);
assign l_31[47]    = ( l_32 [76] & !i[1811]) | ( l_32 [77] &  i[1811]);
assign l_31[48]    = ( l_32 [78] & !i[1811]) | ( l_32 [79] &  i[1811]);
assign l_31[49]    = ( l_32 [80] & !i[1811]) | ( l_32 [81] &  i[1811]);
assign l_31[50]    = ( l_32 [82] & !i[1811]) | ( l_32 [83] &  i[1811]);
assign l_31[51]    = ( l_32 [84] & !i[1811]) | ( l_32 [85] &  i[1811]);
assign l_31[52]    = ( l_32 [86] & !i[1811]) | ( l_32 [87] &  i[1811]);
assign l_31[53]    = ( l_32 [88] & !i[1811]) | ( l_32 [89] &  i[1811]);
assign l_31[54]    = ( l_32 [90] & !i[1811]) | ( l_32 [91] &  i[1811]);
assign l_31[55]    = ( l_32 [92] & !i[1811]) | ( l_32 [93] &  i[1811]);
assign l_31[56]    = ( l_32 [94] & !i[1811]) | ( l_32 [95] &  i[1811]);
assign l_31[57]    = ( l_32 [96] & !i[1811]) | ( l_32 [97] &  i[1811]);
assign l_31[58]    = ( l_32 [98] & !i[1811]) | ( l_32 [99] &  i[1811]);
assign l_31[59]    = ( l_32 [100] & !i[1811]) | ( l_32 [101] &  i[1811]);
assign l_31[60]    = ( l_32 [102] & !i[1811]) | ( l_32 [103] &  i[1811]);
assign l_31[61]    = ( l_32 [104] & !i[1811]) | ( l_32 [105] &  i[1811]);
assign l_31[62]    = ( l_32 [106] & !i[1811]) | ( l_32 [107] &  i[1811]);
assign l_31[63]    = ( l_32 [108] & !i[1811]) | ( l_32 [109] &  i[1811]);
assign l_31[64]    = ( l_32 [110] & !i[1811]) | ( l_32 [111] &  i[1811]);
assign l_31[65]    = ( l_32 [112] & !i[1811]) | ( l_32 [113] &  i[1811]);
assign l_31[66]    = ( l_32 [114] & !i[1811]) | ( l_32 [115] &  i[1811]);
assign l_31[67]    = ( l_32 [116] & !i[1811]) | ( l_32 [117] &  i[1811]);
assign l_31[68]    = ( l_32 [118] & !i[1811]) | ( l_32 [119] &  i[1811]);
assign l_31[69]    = ( l_32 [120] & !i[1811]) | ( l_32 [121] &  i[1811]);
assign l_31[70]    = ( l_32 [122] & !i[1811]) | ( l_32 [123] &  i[1811]);
assign l_31[71]    = ( l_32 [124] & !i[1811]) | ( l_32 [125] &  i[1811]);
assign l_31[72]    = ( l_32 [126] & !i[1811]) | ( l_32 [127] &  i[1811]);
assign l_31[73]    = ( l_32 [128] & !i[1811]) | ( l_32 [129] &  i[1811]);
assign l_31[74]    = ( l_32 [130] & !i[1811]) | ( l_32 [131] &  i[1811]);
assign l_31[75]    = ( l_32 [132] & !i[1811]) | ( l_32 [133] &  i[1811]);
assign l_31[76]    = ( l_32 [134] & !i[1811]) | ( l_32 [135] &  i[1811]);
assign l_31[77]    = ( l_32 [136] & !i[1811]) | ( l_32 [137] &  i[1811]);
assign l_31[78]    = ( l_32 [138] & !i[1811]) | ( l_32 [139] &  i[1811]);
assign l_31[79]    = ( l_32 [140] & !i[1811]) | ( l_32 [141] &  i[1811]);
assign l_31[80]    = ( l_32 [142] & !i[1811]) | ( l_32 [143] &  i[1811]);
assign l_31[81]    = ( l_32 [144] & !i[1811]) | ( l_32 [145] &  i[1811]);
assign l_31[82]    = ( l_32 [146]);
assign l_31[83]    = ( l_32 [147]);
assign l_31[84]    = ( l_32 [148]);
assign l_31[85]    = ( l_32 [149]);
assign l_31[86]    = ( l_32 [150]);
assign l_31[87]    = ( l_32 [151]);
assign l_31[88]    = ( l_32 [152]);
assign l_31[89]    = ( l_32 [153]);
assign l_31[90]    = ( l_32 [154]);
assign l_31[91]    = ( l_32 [155]);
assign l_31[92]    = ( l_32 [156]);
assign l_31[93]    = ( l_32 [157]);
assign l_31[94]    = ( l_32 [158]);
assign l_31[95]    = ( l_32 [159]);
assign l_31[96]    = ( l_32 [160]);
assign l_31[97]    = ( l_32 [161]);
assign l_31[98]    = ( l_32 [162]);
assign l_31[99]    = ( l_32 [163]);
assign l_31[100]    = ( l_32 [164]);
assign l_31[101]    = ( l_32 [165]);
assign l_31[102]    = ( l_32 [166]);
assign l_31[103]    = ( l_32 [167]);
assign l_31[104]    = ( l_32 [168]);
assign l_31[105]    = ( l_32 [169]);
assign l_31[106]    = ( l_32 [170]);
assign l_31[107]    = ( l_32 [171]);
assign l_31[108]    = ( l_32 [172]);
assign l_31[109]    = ( l_32 [173]);
assign l_31[110]    = ( l_32 [174]);
assign l_31[111]    = ( l_32 [175]);
assign l_31[112]    = ( l_32 [176]);
assign l_31[113]    = ( l_32 [177]);
assign l_31[114]    = ( l_32 [178]);
assign l_31[115]    = ( l_32 [179]);
assign l_31[116]    = ( l_32 [180]);
assign l_31[117]    = ( l_32 [181]);
assign l_31[118]    = ( l_32 [182]);
assign l_31[119]    = ( l_32 [183]);
assign l_31[120]    = ( l_32 [184]);
assign l_31[121]    = ( l_32 [185]);
assign l_31[122]    = ( l_32 [186]);
assign l_31[123]    = ( l_32 [187]);
assign l_31[124]    = ( l_32 [188]);
assign l_31[125]    = ( l_32 [189]);
assign l_31[126]    = ( l_32 [190]);
assign l_31[127]    = ( l_32 [191]);
assign l_31[128]    = ( l_32 [192]);
assign l_31[129]    = ( l_32 [193]);
assign l_31[130]    = ( l_32 [194]);
assign l_31[131]    = ( l_32 [195]);
assign l_31[132]    = ( l_32 [196]);
assign l_31[133]    = ( l_32 [197]);
assign l_31[134]    = ( l_32 [198]);
assign l_31[135]    = ( l_32 [199]);
assign l_31[136]    = ( l_32 [200]);
assign l_31[137]    = ( l_32 [201]);
assign l_31[138]    = ( l_32 [202]);
assign l_31[139]    = ( l_32 [203]);
assign l_31[140]    = ( l_32 [204]);
assign l_31[141]    = ( l_32 [205]);
assign l_31[142]    = ( l_32 [206]);
assign l_31[143]    = ( l_32 [207]);
assign l_31[144]    = ( l_32 [208]);
assign l_31[145]    = ( l_32 [209]);
assign l_31[146]    = ( l_32 [210]);
assign l_31[147]    = ( l_32 [211]);
assign l_31[148]    = ( l_32 [212]);
assign l_31[149]    = ( l_32 [213]);
assign l_31[150]    = ( l_32 [214]);
assign l_31[151]    = ( l_32 [215]);
assign l_31[152]    = ( l_32 [216]);
assign l_31[153]    = ( l_32 [217]);
assign l_31[154]    = ( l_32 [218]);
assign l_31[155]    = ( l_32 [219]);
assign l_31[156]    = ( l_32 [220]);
assign l_31[157]    = ( l_32 [221]);
assign l_31[158]    = ( l_32 [222]);
assign l_31[159]    = ( l_32 [223]);
assign l_31[160]    = ( l_32 [224]);
assign l_31[161]    = ( l_32 [225]);
assign l_31[162]    = ( l_32 [226]);
assign l_31[163]    = ( l_32 [227]);
assign l_31[164]    = ( l_32 [228]);
assign l_31[165]    = ( l_32 [229]);
assign l_31[166]    = ( l_32 [230]);
assign l_31[167]    = ( l_32 [231]);
assign l_31[168]    = ( l_32 [232]);
assign l_31[169]    = ( l_32 [233]);
assign l_31[170]    = ( l_32 [234]);
assign l_31[171]    = ( l_32 [235]);
assign l_31[172]    = ( l_32 [236]);
assign l_31[173]    = ( l_32 [237]);
assign l_31[174]    = ( l_32 [238]);
assign l_31[175]    = ( l_32 [239]);
assign l_31[176]    = ( l_32 [240]);
assign l_31[177]    = ( l_32 [241]);
assign l_31[178]    = ( l_32 [242]);
assign l_31[179]    = ( l_32 [243]);
assign l_31[180]    = ( l_32 [244]);
assign l_31[181]    = ( l_32 [245]);
assign l_31[182]    = ( l_32 [246]);
assign l_31[183]    = ( l_32 [247]);
assign l_31[184]    = ( l_32 [248]);
assign l_31[185]    = ( l_32 [249]);
assign l_31[186]    = ( l_32 [250]);
assign l_31[187]    = ( l_32 [251]);
assign l_31[188]    = ( l_32 [252]);
assign l_31[189]    = ( l_32 [253]);
assign l_31[190]    = ( l_32 [254]);
assign l_31[191]    = ( l_32 [255]);
assign l_31[192]    = ( l_32 [256]);
assign l_31[193]    = ( l_32 [257]);
assign l_31[194]    = ( l_32 [258]);
assign l_31[195]    = ( l_32 [259]);
assign l_31[196]    = ( l_32 [260]);
assign l_31[197]    = ( l_32 [261]);
assign l_31[198]    = ( l_32 [262]);
assign l_31[199]    = ( l_32 [263]);
assign l_31[200]    = ( l_32 [264]);
assign l_31[201]    = ( l_32 [265]);
assign l_31[202]    = ( l_32 [266]);
assign l_31[203]    = ( l_32 [267]);
assign l_31[204]    = ( l_32 [268]);
assign l_31[205]    = ( l_32 [269]);
assign l_31[206]    = ( l_32 [270]);
assign l_31[207]    = ( l_32 [271]);
assign l_31[208]    = ( l_32 [272]);
assign l_31[209]    = ( l_32 [273]);
assign l_32[0]    = ( l_33 [0]);
assign l_32[1]    = ( l_33 [1] & !i[1807]);
assign l_32[2]    = ( l_33 [2] & !i[1807]);
assign l_32[3]    = (!i[1807]) | ( l_33 [3] &  i[1807]);
assign l_32[4]    = (!i[1807]) | ( l_33 [4] &  i[1807]);
assign l_32[5]    = ( l_33 [5] & !i[1807]);
assign l_32[6]    = ( l_33 [6] & !i[1807]);
assign l_32[7]    = (!i[1807]) | ( l_33 [7] &  i[1807]);
assign l_32[8]    = (!i[1807]) | ( l_33 [8] &  i[1807]);
assign l_32[9]    = ( l_33 [9] & !i[1807]) | ( l_33 [10] &  i[1807]);
assign l_32[10]    = ( l_33 [10]);
assign l_32[11]    = ( l_33 [11] & !i[1807]) | ( l_33 [10] &  i[1807]);
assign l_32[12]    = ( l_33 [10] & !i[1807]) | ( l_33 [12] &  i[1807]);
assign l_32[13]    = ( l_33 [10] & !i[1807]) | ( l_33 [13] &  i[1807]);
assign l_32[14]    = ( l_33 [14] & !i[1807]) | ( l_33 [10] &  i[1807]);
assign l_32[15]    = ( l_33 [15] & !i[1807]) | ( l_33 [10] &  i[1807]);
assign l_32[16]    = ( l_33 [10] & !i[1807]) | ( l_33 [16] &  i[1807]);
assign l_32[17]    = ( l_33 [10] & !i[1807]) | ( l_33 [17] &  i[1807]);
assign l_32[18]    = ( l_33 [18] & !i[1807]) | ( l_33 [19] &  i[1807]);
assign l_32[19]    = ( l_33 [20] & !i[1807]) | ( l_33 [21] &  i[1807]);
assign l_32[20]    = ( l_33 [22] & !i[1807]) | ( l_33 [23] &  i[1807]);
assign l_32[21]    = ( l_33 [24] & !i[1807]) | ( l_33 [25] &  i[1807]);
assign l_32[22]    = ( l_33 [26] & !i[1807]) | ( l_33 [27] &  i[1807]);
assign l_32[23]    = ( l_33 [28] & !i[1807]) | ( l_33 [29] &  i[1807]);
assign l_32[24]    = ( l_33 [30] & !i[1807]) | ( l_33 [31] &  i[1807]);
assign l_32[25]    = ( l_33 [32] & !i[1807]) | ( l_33 [33] &  i[1807]);
assign l_32[26]    = ( l_33 [34] & !i[1807]) | ( l_33 [35] &  i[1807]);
assign l_32[27]    = ( l_33 [36] & !i[1807]) | ( l_33 [37] &  i[1807]);
assign l_32[28]    = ( l_33 [38] & !i[1807]) | ( l_33 [39] &  i[1807]);
assign l_32[29]    = ( l_33 [40] & !i[1807]) | ( l_33 [41] &  i[1807]);
assign l_32[30]    = ( l_33 [42] & !i[1807]) | ( l_33 [43] &  i[1807]);
assign l_32[31]    = ( l_33 [44] & !i[1807]) | ( l_33 [45] &  i[1807]);
assign l_32[32]    = ( l_33 [46] & !i[1807]) | ( l_33 [47] &  i[1807]);
assign l_32[33]    = ( l_33 [48] & !i[1807]) | ( l_33 [49] &  i[1807]);
assign l_32[34]    = ( l_33 [50] & !i[1807]) | ( l_33 [51] &  i[1807]);
assign l_32[35]    = ( l_33 [52] & !i[1807]) | ( l_33 [53] &  i[1807]);
assign l_32[36]    = ( l_33 [54] & !i[1807]) | ( l_33 [55] &  i[1807]);
assign l_32[37]    = ( l_33 [56] & !i[1807]) | ( l_33 [57] &  i[1807]);
assign l_32[38]    = ( l_33 [58] & !i[1807]) | ( l_33 [59] &  i[1807]);
assign l_32[39]    = ( l_33 [60] & !i[1807]) | ( l_33 [61] &  i[1807]);
assign l_32[40]    = ( l_33 [62] & !i[1807]) | ( l_33 [63] &  i[1807]);
assign l_32[41]    = ( l_33 [64] & !i[1807]) | ( l_33 [65] &  i[1807]);
assign l_32[42]    = ( l_33 [66] & !i[1807]) | ( l_33 [67] &  i[1807]);
assign l_32[43]    = ( l_33 [68] & !i[1807]) | ( l_33 [69] &  i[1807]);
assign l_32[44]    = ( l_33 [70] & !i[1807]) | ( l_33 [71] &  i[1807]);
assign l_32[45]    = ( l_33 [72] & !i[1807]) | ( l_33 [73] &  i[1807]);
assign l_32[46]    = ( l_33 [74] & !i[1807]) | ( l_33 [75] &  i[1807]);
assign l_32[47]    = ( l_33 [76] & !i[1807]) | ( l_33 [77] &  i[1807]);
assign l_32[48]    = ( l_33 [78] & !i[1807]) | ( l_33 [79] &  i[1807]);
assign l_32[49]    = ( l_33 [80] & !i[1807]) | ( l_33 [81] &  i[1807]);
assign l_32[50]    = ( l_33 [82] & !i[1807]) | ( l_33 [83] &  i[1807]);
assign l_32[51]    = ( l_33 [84] & !i[1807]) | ( l_33 [85] &  i[1807]);
assign l_32[52]    = ( l_33 [86] & !i[1807]) | ( l_33 [87] &  i[1807]);
assign l_32[53]    = ( l_33 [88] & !i[1807]) | ( l_33 [89] &  i[1807]);
assign l_32[54]    = ( l_33 [90] & !i[1807]) | ( l_33 [91] &  i[1807]);
assign l_32[55]    = ( l_33 [92] & !i[1807]) | ( l_33 [93] &  i[1807]);
assign l_32[56]    = ( l_33 [94] & !i[1807]) | ( l_33 [95] &  i[1807]);
assign l_32[57]    = ( l_33 [96] & !i[1807]) | ( l_33 [97] &  i[1807]);
assign l_32[58]    = ( l_33 [98] & !i[1807]) | ( l_33 [99] &  i[1807]);
assign l_32[59]    = ( l_33 [100] & !i[1807]) | ( l_33 [101] &  i[1807]);
assign l_32[60]    = ( l_33 [102] & !i[1807]) | ( l_33 [103] &  i[1807]);
assign l_32[61]    = ( l_33 [104] & !i[1807]) | ( l_33 [105] &  i[1807]);
assign l_32[62]    = ( l_33 [106] & !i[1807]) | ( l_33 [107] &  i[1807]);
assign l_32[63]    = ( l_33 [108] & !i[1807]) | ( l_33 [109] &  i[1807]);
assign l_32[64]    = ( l_33 [110] & !i[1807]) | ( l_33 [111] &  i[1807]);
assign l_32[65]    = ( l_33 [112] & !i[1807]) | ( l_33 [113] &  i[1807]);
assign l_32[66]    = ( l_33 [114] & !i[1807]) | ( l_33 [115] &  i[1807]);
assign l_32[67]    = ( l_33 [116] & !i[1807]) | ( l_33 [117] &  i[1807]);
assign l_32[68]    = ( l_33 [118] & !i[1807]) | ( l_33 [119] &  i[1807]);
assign l_32[69]    = ( l_33 [120] & !i[1807]) | ( l_33 [121] &  i[1807]);
assign l_32[70]    = ( l_33 [122] & !i[1807]) | ( l_33 [123] &  i[1807]);
assign l_32[71]    = ( l_33 [124] & !i[1807]) | ( l_33 [125] &  i[1807]);
assign l_32[72]    = ( l_33 [126] & !i[1807]) | ( l_33 [127] &  i[1807]);
assign l_32[73]    = ( l_33 [128] & !i[1807]) | ( l_33 [129] &  i[1807]);
assign l_32[74]    = ( l_33 [130] & !i[1807]) | ( l_33 [131] &  i[1807]);
assign l_32[75]    = ( l_33 [132] & !i[1807]) | ( l_33 [133] &  i[1807]);
assign l_32[76]    = ( l_33 [134] & !i[1807]) | ( l_33 [135] &  i[1807]);
assign l_32[77]    = ( l_33 [136] & !i[1807]) | ( l_33 [137] &  i[1807]);
assign l_32[78]    = ( l_33 [138] & !i[1807]) | ( l_33 [139] &  i[1807]);
assign l_32[79]    = ( l_33 [140] & !i[1807]) | ( l_33 [141] &  i[1807]);
assign l_32[80]    = ( l_33 [142] & !i[1807]) | ( l_33 [143] &  i[1807]);
assign l_32[81]    = ( l_33 [144] & !i[1807]) | ( l_33 [145] &  i[1807]);
assign l_32[82]    = ( l_33 [146] & !i[1807]) | ( l_33 [147] &  i[1807]);
assign l_32[83]    = ( l_33 [148] & !i[1807]) | ( l_33 [149] &  i[1807]);
assign l_32[84]    = ( l_33 [150] & !i[1807]) | ( l_33 [151] &  i[1807]);
assign l_32[85]    = ( l_33 [152] & !i[1807]) | ( l_33 [153] &  i[1807]);
assign l_32[86]    = ( l_33 [154] & !i[1807]) | ( l_33 [155] &  i[1807]);
assign l_32[87]    = ( l_33 [156] & !i[1807]) | ( l_33 [157] &  i[1807]);
assign l_32[88]    = ( l_33 [158] & !i[1807]) | ( l_33 [159] &  i[1807]);
assign l_32[89]    = ( l_33 [160] & !i[1807]) | ( l_33 [161] &  i[1807]);
assign l_32[90]    = ( l_33 [162] & !i[1807]) | ( l_33 [163] &  i[1807]);
assign l_32[91]    = ( l_33 [164] & !i[1807]) | ( l_33 [165] &  i[1807]);
assign l_32[92]    = ( l_33 [166] & !i[1807]) | ( l_33 [167] &  i[1807]);
assign l_32[93]    = ( l_33 [168] & !i[1807]) | ( l_33 [169] &  i[1807]);
assign l_32[94]    = ( l_33 [170] & !i[1807]) | ( l_33 [171] &  i[1807]);
assign l_32[95]    = ( l_33 [172] & !i[1807]) | ( l_33 [173] &  i[1807]);
assign l_32[96]    = ( l_33 [174] & !i[1807]) | ( l_33 [175] &  i[1807]);
assign l_32[97]    = ( l_33 [176] & !i[1807]) | ( l_33 [177] &  i[1807]);
assign l_32[98]    = ( l_33 [178] & !i[1807]) | ( l_33 [179] &  i[1807]);
assign l_32[99]    = ( l_33 [180] & !i[1807]) | ( l_33 [181] &  i[1807]);
assign l_32[100]    = ( l_33 [182] & !i[1807]) | ( l_33 [183] &  i[1807]);
assign l_32[101]    = ( l_33 [184] & !i[1807]) | ( l_33 [185] &  i[1807]);
assign l_32[102]    = ( l_33 [186] & !i[1807]) | ( l_33 [187] &  i[1807]);
assign l_32[103]    = ( l_33 [188] & !i[1807]) | ( l_33 [189] &  i[1807]);
assign l_32[104]    = ( l_33 [190] & !i[1807]) | ( l_33 [191] &  i[1807]);
assign l_32[105]    = ( l_33 [192] & !i[1807]) | ( l_33 [193] &  i[1807]);
assign l_32[106]    = ( l_33 [194] & !i[1807]) | ( l_33 [195] &  i[1807]);
assign l_32[107]    = ( l_33 [196] & !i[1807]) | ( l_33 [197] &  i[1807]);
assign l_32[108]    = ( l_33 [198] & !i[1807]) | ( l_33 [199] &  i[1807]);
assign l_32[109]    = ( l_33 [200] & !i[1807]) | ( l_33 [201] &  i[1807]);
assign l_32[110]    = ( l_33 [202] & !i[1807]) | ( l_33 [203] &  i[1807]);
assign l_32[111]    = ( l_33 [204] & !i[1807]) | ( l_33 [205] &  i[1807]);
assign l_32[112]    = ( l_33 [206] & !i[1807]) | ( l_33 [207] &  i[1807]);
assign l_32[113]    = ( l_33 [208] & !i[1807]) | ( l_33 [209] &  i[1807]);
assign l_32[114]    = ( l_33 [210] & !i[1807]) | ( l_33 [211] &  i[1807]);
assign l_32[115]    = ( l_33 [212] & !i[1807]) | ( l_33 [213] &  i[1807]);
assign l_32[116]    = ( l_33 [214] & !i[1807]) | ( l_33 [215] &  i[1807]);
assign l_32[117]    = ( l_33 [216] & !i[1807]) | ( l_33 [217] &  i[1807]);
assign l_32[118]    = ( l_33 [218] & !i[1807]) | ( l_33 [219] &  i[1807]);
assign l_32[119]    = ( l_33 [220] & !i[1807]) | ( l_33 [221] &  i[1807]);
assign l_32[120]    = ( l_33 [222] & !i[1807]) | ( l_33 [223] &  i[1807]);
assign l_32[121]    = ( l_33 [224] & !i[1807]) | ( l_33 [225] &  i[1807]);
assign l_32[122]    = ( l_33 [226] & !i[1807]) | ( l_33 [227] &  i[1807]);
assign l_32[123]    = ( l_33 [228] & !i[1807]) | ( l_33 [229] &  i[1807]);
assign l_32[124]    = ( l_33 [230] & !i[1807]) | ( l_33 [231] &  i[1807]);
assign l_32[125]    = ( l_33 [232] & !i[1807]) | ( l_33 [233] &  i[1807]);
assign l_32[126]    = ( l_33 [234] & !i[1807]) | ( l_33 [235] &  i[1807]);
assign l_32[127]    = ( l_33 [236] & !i[1807]) | ( l_33 [237] &  i[1807]);
assign l_32[128]    = ( l_33 [238] & !i[1807]) | ( l_33 [239] &  i[1807]);
assign l_32[129]    = ( l_33 [240] & !i[1807]) | ( l_33 [241] &  i[1807]);
assign l_32[130]    = ( l_33 [242] & !i[1807]) | ( l_33 [243] &  i[1807]);
assign l_32[131]    = ( l_33 [244] & !i[1807]) | ( l_33 [245] &  i[1807]);
assign l_32[132]    = ( l_33 [246] & !i[1807]) | ( l_33 [247] &  i[1807]);
assign l_32[133]    = ( l_33 [248] & !i[1807]) | ( l_33 [249] &  i[1807]);
assign l_32[134]    = ( l_33 [250] & !i[1807]) | ( l_33 [251] &  i[1807]);
assign l_32[135]    = ( l_33 [252] & !i[1807]) | ( l_33 [253] &  i[1807]);
assign l_32[136]    = ( l_33 [254] & !i[1807]) | ( l_33 [255] &  i[1807]);
assign l_32[137]    = ( l_33 [256] & !i[1807]) | ( l_33 [257] &  i[1807]);
assign l_32[138]    = ( l_33 [258] & !i[1807]) | ( l_33 [259] &  i[1807]);
assign l_32[139]    = ( l_33 [260] & !i[1807]) | ( l_33 [261] &  i[1807]);
assign l_32[140]    = ( l_33 [262] & !i[1807]) | ( l_33 [263] &  i[1807]);
assign l_32[141]    = ( l_33 [264] & !i[1807]) | ( l_33 [265] &  i[1807]);
assign l_32[142]    = ( l_33 [266] & !i[1807]) | ( l_33 [267] &  i[1807]);
assign l_32[143]    = ( l_33 [268] & !i[1807]) | ( l_33 [269] &  i[1807]);
assign l_32[144]    = ( l_33 [270] & !i[1807]) | ( l_33 [271] &  i[1807]);
assign l_32[145]    = ( l_33 [272] & !i[1807]) | ( l_33 [273] &  i[1807]);
assign l_32[146]    = ( l_33 [274]);
assign l_32[147]    = ( l_33 [275]);
assign l_32[148]    = ( l_33 [276]);
assign l_32[149]    = ( l_33 [277]);
assign l_32[150]    = ( l_33 [278]);
assign l_32[151]    = ( l_33 [279]);
assign l_32[152]    = ( l_33 [280]);
assign l_32[153]    = ( l_33 [281]);
assign l_32[154]    = ( l_33 [282]);
assign l_32[155]    = ( l_33 [283]);
assign l_32[156]    = ( l_33 [284]);
assign l_32[157]    = ( l_33 [285]);
assign l_32[158]    = ( l_33 [286]);
assign l_32[159]    = ( l_33 [287]);
assign l_32[160]    = ( l_33 [288]);
assign l_32[161]    = ( l_33 [289]);
assign l_32[162]    = ( l_33 [290]);
assign l_32[163]    = ( l_33 [291]);
assign l_32[164]    = ( l_33 [292]);
assign l_32[165]    = ( l_33 [293]);
assign l_32[166]    = ( l_33 [294]);
assign l_32[167]    = ( l_33 [295]);
assign l_32[168]    = ( l_33 [296]);
assign l_32[169]    = ( l_33 [297]);
assign l_32[170]    = ( l_33 [298]);
assign l_32[171]    = ( l_33 [299]);
assign l_32[172]    = ( l_33 [300]);
assign l_32[173]    = ( l_33 [301]);
assign l_32[174]    = ( l_33 [302]);
assign l_32[175]    = ( l_33 [303]);
assign l_32[176]    = ( l_33 [304]);
assign l_32[177]    = ( l_33 [305]);
assign l_32[178]    = ( l_33 [306]);
assign l_32[179]    = ( l_33 [307]);
assign l_32[180]    = ( l_33 [308]);
assign l_32[181]    = ( l_33 [309]);
assign l_32[182]    = ( l_33 [310]);
assign l_32[183]    = ( l_33 [311]);
assign l_32[184]    = ( l_33 [312]);
assign l_32[185]    = ( l_33 [313]);
assign l_32[186]    = ( l_33 [314]);
assign l_32[187]    = ( l_33 [315]);
assign l_32[188]    = ( l_33 [316]);
assign l_32[189]    = ( l_33 [317]);
assign l_32[190]    = ( l_33 [318]);
assign l_32[191]    = ( l_33 [319]);
assign l_32[192]    = ( l_33 [320]);
assign l_32[193]    = ( l_33 [321]);
assign l_32[194]    = ( l_33 [322]);
assign l_32[195]    = ( l_33 [323]);
assign l_32[196]    = ( l_33 [324]);
assign l_32[197]    = ( l_33 [325]);
assign l_32[198]    = ( l_33 [326]);
assign l_32[199]    = ( l_33 [327]);
assign l_32[200]    = ( l_33 [328]);
assign l_32[201]    = ( l_33 [329]);
assign l_32[202]    = ( l_33 [330]);
assign l_32[203]    = ( l_33 [331]);
assign l_32[204]    = ( l_33 [332]);
assign l_32[205]    = ( l_33 [333]);
assign l_32[206]    = ( l_33 [334]);
assign l_32[207]    = ( l_33 [335]);
assign l_32[208]    = ( l_33 [336]);
assign l_32[209]    = ( l_33 [337]);
assign l_32[210]    = ( l_33 [338]);
assign l_32[211]    = ( l_33 [339]);
assign l_32[212]    = ( l_33 [340]);
assign l_32[213]    = ( l_33 [341]);
assign l_32[214]    = ( l_33 [342]);
assign l_32[215]    = ( l_33 [343]);
assign l_32[216]    = ( l_33 [344]);
assign l_32[217]    = ( l_33 [345]);
assign l_32[218]    = ( l_33 [346]);
assign l_32[219]    = ( l_33 [347]);
assign l_32[220]    = ( l_33 [348]);
assign l_32[221]    = ( l_33 [349]);
assign l_32[222]    = ( l_33 [350]);
assign l_32[223]    = ( l_33 [351]);
assign l_32[224]    = ( l_33 [352]);
assign l_32[225]    = ( l_33 [353]);
assign l_32[226]    = ( l_33 [354]);
assign l_32[227]    = ( l_33 [355]);
assign l_32[228]    = ( l_33 [356]);
assign l_32[229]    = ( l_33 [357]);
assign l_32[230]    = ( l_33 [358]);
assign l_32[231]    = ( l_33 [359]);
assign l_32[232]    = ( l_33 [360]);
assign l_32[233]    = ( l_33 [361]);
assign l_32[234]    = ( l_33 [362]);
assign l_32[235]    = ( l_33 [363]);
assign l_32[236]    = ( l_33 [364]);
assign l_32[237]    = ( l_33 [365]);
assign l_32[238]    = ( l_33 [366]);
assign l_32[239]    = ( l_33 [367]);
assign l_32[240]    = ( l_33 [368]);
assign l_32[241]    = ( l_33 [369]);
assign l_32[242]    = ( l_33 [370]);
assign l_32[243]    = ( l_33 [371]);
assign l_32[244]    = ( l_33 [372]);
assign l_32[245]    = ( l_33 [373]);
assign l_32[246]    = ( l_33 [374]);
assign l_32[247]    = ( l_33 [375]);
assign l_32[248]    = ( l_33 [376]);
assign l_32[249]    = ( l_33 [377]);
assign l_32[250]    = ( l_33 [378]);
assign l_32[251]    = ( l_33 [379]);
assign l_32[252]    = ( l_33 [380]);
assign l_32[253]    = ( l_33 [381]);
assign l_32[254]    = ( l_33 [382]);
assign l_32[255]    = ( l_33 [383]);
assign l_32[256]    = ( l_33 [384]);
assign l_32[257]    = ( l_33 [385]);
assign l_32[258]    = ( l_33 [386]);
assign l_32[259]    = ( l_33 [387]);
assign l_32[260]    = ( l_33 [388]);
assign l_32[261]    = ( l_33 [389]);
assign l_32[262]    = ( l_33 [390]);
assign l_32[263]    = ( l_33 [391]);
assign l_32[264]    = ( l_33 [392]);
assign l_32[265]    = ( l_33 [393]);
assign l_32[266]    = ( l_33 [394]);
assign l_32[267]    = ( l_33 [395]);
assign l_32[268]    = ( l_33 [396]);
assign l_32[269]    = ( l_33 [397]);
assign l_32[270]    = ( l_33 [398]);
assign l_32[271]    = ( l_33 [399]);
assign l_32[272]    = ( l_33 [400]);
assign l_32[273]    = ( l_33 [401]);
assign l_33[0]    = ( l_34 [0]);
assign l_33[1]    = ( l_34 [1] & !i[1818]);
assign l_33[2]    = ( l_34 [2] & !i[1818]);
assign l_33[3]    = (!i[1818]) | ( l_34 [3] &  i[1818]);
assign l_33[4]    = (!i[1818]) | ( l_34 [4] &  i[1818]);
assign l_33[5]    = ( l_34 [5] & !i[1818]);
assign l_33[6]    = ( l_34 [6] & !i[1818]);
assign l_33[7]    = (!i[1818]) | ( l_34 [7] &  i[1818]);
assign l_33[8]    = (!i[1818]) | ( l_34 [8] &  i[1818]);
assign l_33[9]    = ( l_34 [9] & !i[1818]) | ( l_34 [10] &  i[1818]);
assign l_33[10]    = ( l_34 [10]);
assign l_33[11]    = ( l_34 [11] & !i[1818]) | ( l_34 [10] &  i[1818]);
assign l_33[12]    = ( l_34 [10] & !i[1818]) | ( l_34 [12] &  i[1818]);
assign l_33[13]    = ( l_34 [10] & !i[1818]) | ( l_34 [13] &  i[1818]);
assign l_33[14]    = ( l_34 [14] & !i[1818]) | ( l_34 [10] &  i[1818]);
assign l_33[15]    = ( l_34 [15] & !i[1818]) | ( l_34 [10] &  i[1818]);
assign l_33[16]    = ( l_34 [10] & !i[1818]) | ( l_34 [16] &  i[1818]);
assign l_33[17]    = ( l_34 [10] & !i[1818]) | ( l_34 [17] &  i[1818]);
assign l_33[18]    = ( l_34 [18]);
assign l_33[19]    = ( l_34 [19]);
assign l_33[20]    = ( l_34 [20]);
assign l_33[21]    = ( l_34 [21]);
assign l_33[22]    = ( l_34 [22]);
assign l_33[23]    = ( l_34 [23]);
assign l_33[24]    = ( l_34 [24]);
assign l_33[25]    = ( l_34 [25]);
assign l_33[26]    = ( l_34 [26]);
assign l_33[27]    = ( l_34 [27]);
assign l_33[28]    = ( l_34 [28]);
assign l_33[29]    = ( l_34 [29]);
assign l_33[30]    = ( l_34 [30]);
assign l_33[31]    = ( l_34 [31]);
assign l_33[32]    = ( l_34 [32]);
assign l_33[33]    = ( l_34 [33]);
assign l_33[34]    = ( l_34 [34]);
assign l_33[35]    = ( l_34 [35]);
assign l_33[36]    = ( l_34 [36]);
assign l_33[37]    = ( l_34 [37]);
assign l_33[38]    = ( l_34 [38]);
assign l_33[39]    = ( l_34 [39]);
assign l_33[40]    = ( l_34 [40]);
assign l_33[41]    = ( l_34 [41]);
assign l_33[42]    = ( l_34 [42]);
assign l_33[43]    = ( l_34 [43]);
assign l_33[44]    = ( l_34 [44]);
assign l_33[45]    = ( l_34 [45]);
assign l_33[46]    = ( l_34 [46]);
assign l_33[47]    = ( l_34 [47]);
assign l_33[48]    = ( l_34 [48]);
assign l_33[49]    = ( l_34 [49]);
assign l_33[50]    = ( l_34 [50]);
assign l_33[51]    = ( l_34 [51]);
assign l_33[52]    = ( l_34 [52]);
assign l_33[53]    = ( l_34 [53]);
assign l_33[54]    = ( l_34 [54]);
assign l_33[55]    = ( l_34 [55]);
assign l_33[56]    = ( l_34 [56]);
assign l_33[57]    = ( l_34 [57]);
assign l_33[58]    = ( l_34 [58]);
assign l_33[59]    = ( l_34 [59]);
assign l_33[60]    = ( l_34 [60]);
assign l_33[61]    = ( l_34 [61]);
assign l_33[62]    = ( l_34 [62]);
assign l_33[63]    = ( l_34 [63]);
assign l_33[64]    = ( l_34 [64]);
assign l_33[65]    = ( l_34 [65]);
assign l_33[66]    = ( l_34 [66]);
assign l_33[67]    = ( l_34 [67]);
assign l_33[68]    = ( l_34 [68]);
assign l_33[69]    = ( l_34 [69]);
assign l_33[70]    = ( l_34 [70]);
assign l_33[71]    = ( l_34 [71]);
assign l_33[72]    = ( l_34 [72]);
assign l_33[73]    = ( l_34 [73]);
assign l_33[74]    = ( l_34 [74]);
assign l_33[75]    = ( l_34 [75]);
assign l_33[76]    = ( l_34 [76]);
assign l_33[77]    = ( l_34 [77]);
assign l_33[78]    = ( l_34 [78]);
assign l_33[79]    = ( l_34 [79]);
assign l_33[80]    = ( l_34 [80]);
assign l_33[81]    = ( l_34 [81]);
assign l_33[82]    = ( l_34 [82]);
assign l_33[83]    = ( l_34 [83]);
assign l_33[84]    = ( l_34 [84]);
assign l_33[85]    = ( l_34 [85]);
assign l_33[86]    = ( l_34 [86]);
assign l_33[87]    = ( l_34 [87]);
assign l_33[88]    = ( l_34 [88]);
assign l_33[89]    = ( l_34 [89]);
assign l_33[90]    = ( l_34 [90]);
assign l_33[91]    = ( l_34 [91]);
assign l_33[92]    = ( l_34 [92]);
assign l_33[93]    = ( l_34 [93]);
assign l_33[94]    = ( l_34 [94]);
assign l_33[95]    = ( l_34 [95]);
assign l_33[96]    = ( l_34 [96]);
assign l_33[97]    = ( l_34 [97]);
assign l_33[98]    = ( l_34 [98]);
assign l_33[99]    = ( l_34 [99]);
assign l_33[100]    = ( l_34 [100]);
assign l_33[101]    = ( l_34 [101]);
assign l_33[102]    = ( l_34 [102]);
assign l_33[103]    = ( l_34 [103]);
assign l_33[104]    = ( l_34 [104]);
assign l_33[105]    = ( l_34 [105]);
assign l_33[106]    = ( l_34 [106]);
assign l_33[107]    = ( l_34 [107]);
assign l_33[108]    = ( l_34 [108]);
assign l_33[109]    = ( l_34 [109]);
assign l_33[110]    = ( l_34 [110]);
assign l_33[111]    = ( l_34 [111]);
assign l_33[112]    = ( l_34 [112]);
assign l_33[113]    = ( l_34 [113]);
assign l_33[114]    = ( l_34 [114]);
assign l_33[115]    = ( l_34 [115]);
assign l_33[116]    = ( l_34 [116]);
assign l_33[117]    = ( l_34 [117]);
assign l_33[118]    = ( l_34 [118]);
assign l_33[119]    = ( l_34 [119]);
assign l_33[120]    = ( l_34 [120]);
assign l_33[121]    = ( l_34 [121]);
assign l_33[122]    = ( l_34 [122]);
assign l_33[123]    = ( l_34 [123]);
assign l_33[124]    = ( l_34 [124]);
assign l_33[125]    = ( l_34 [125]);
assign l_33[126]    = ( l_34 [126]);
assign l_33[127]    = ( l_34 [127]);
assign l_33[128]    = ( l_34 [128]);
assign l_33[129]    = ( l_34 [129]);
assign l_33[130]    = ( l_34 [130]);
assign l_33[131]    = ( l_34 [131]);
assign l_33[132]    = ( l_34 [132]);
assign l_33[133]    = ( l_34 [133]);
assign l_33[134]    = ( l_34 [134]);
assign l_33[135]    = ( l_34 [135]);
assign l_33[136]    = ( l_34 [136]);
assign l_33[137]    = ( l_34 [137]);
assign l_33[138]    = ( l_34 [138]);
assign l_33[139]    = ( l_34 [139]);
assign l_33[140]    = ( l_34 [140]);
assign l_33[141]    = ( l_34 [141]);
assign l_33[142]    = ( l_34 [142]);
assign l_33[143]    = ( l_34 [143]);
assign l_33[144]    = ( l_34 [144]);
assign l_33[145]    = ( l_34 [145]);
assign l_33[146]    = ( l_34 [146]);
assign l_33[147]    = ( l_34 [147]);
assign l_33[148]    = ( l_34 [148]);
assign l_33[149]    = ( l_34 [149]);
assign l_33[150]    = ( l_34 [150]);
assign l_33[151]    = ( l_34 [151]);
assign l_33[152]    = ( l_34 [152]);
assign l_33[153]    = ( l_34 [153]);
assign l_33[154]    = ( l_34 [154]);
assign l_33[155]    = ( l_34 [155]);
assign l_33[156]    = ( l_34 [156]);
assign l_33[157]    = ( l_34 [157]);
assign l_33[158]    = ( l_34 [158]);
assign l_33[159]    = ( l_34 [159]);
assign l_33[160]    = ( l_34 [160]);
assign l_33[161]    = ( l_34 [161]);
assign l_33[162]    = ( l_34 [162]);
assign l_33[163]    = ( l_34 [163]);
assign l_33[164]    = ( l_34 [164]);
assign l_33[165]    = ( l_34 [165]);
assign l_33[166]    = ( l_34 [166]);
assign l_33[167]    = ( l_34 [167]);
assign l_33[168]    = ( l_34 [168]);
assign l_33[169]    = ( l_34 [169]);
assign l_33[170]    = ( l_34 [170]);
assign l_33[171]    = ( l_34 [171]);
assign l_33[172]    = ( l_34 [172]);
assign l_33[173]    = ( l_34 [173]);
assign l_33[174]    = ( l_34 [174]);
assign l_33[175]    = ( l_34 [175]);
assign l_33[176]    = ( l_34 [176]);
assign l_33[177]    = ( l_34 [177]);
assign l_33[178]    = ( l_34 [178]);
assign l_33[179]    = ( l_34 [179]);
assign l_33[180]    = ( l_34 [180]);
assign l_33[181]    = ( l_34 [181]);
assign l_33[182]    = ( l_34 [182]);
assign l_33[183]    = ( l_34 [183]);
assign l_33[184]    = ( l_34 [184]);
assign l_33[185]    = ( l_34 [185]);
assign l_33[186]    = ( l_34 [186]);
assign l_33[187]    = ( l_34 [187]);
assign l_33[188]    = ( l_34 [188]);
assign l_33[189]    = ( l_34 [189]);
assign l_33[190]    = ( l_34 [190]);
assign l_33[191]    = ( l_34 [191]);
assign l_33[192]    = ( l_34 [192]);
assign l_33[193]    = ( l_34 [193]);
assign l_33[194]    = ( l_34 [194]);
assign l_33[195]    = ( l_34 [195]);
assign l_33[196]    = ( l_34 [196]);
assign l_33[197]    = ( l_34 [197]);
assign l_33[198]    = ( l_34 [198]);
assign l_33[199]    = ( l_34 [199]);
assign l_33[200]    = ( l_34 [200]);
assign l_33[201]    = ( l_34 [201]);
assign l_33[202]    = ( l_34 [202]);
assign l_33[203]    = ( l_34 [203]);
assign l_33[204]    = ( l_34 [204]);
assign l_33[205]    = ( l_34 [205]);
assign l_33[206]    = ( l_34 [206]);
assign l_33[207]    = ( l_34 [207]);
assign l_33[208]    = ( l_34 [208]);
assign l_33[209]    = ( l_34 [209]);
assign l_33[210]    = ( l_34 [210]);
assign l_33[211]    = ( l_34 [211]);
assign l_33[212]    = ( l_34 [212]);
assign l_33[213]    = ( l_34 [213]);
assign l_33[214]    = ( l_34 [214]);
assign l_33[215]    = ( l_34 [215]);
assign l_33[216]    = ( l_34 [216]);
assign l_33[217]    = ( l_34 [217]);
assign l_33[218]    = ( l_34 [218]);
assign l_33[219]    = ( l_34 [219]);
assign l_33[220]    = ( l_34 [220]);
assign l_33[221]    = ( l_34 [221]);
assign l_33[222]    = ( l_34 [222]);
assign l_33[223]    = ( l_34 [223]);
assign l_33[224]    = ( l_34 [224]);
assign l_33[225]    = ( l_34 [225]);
assign l_33[226]    = ( l_34 [226]);
assign l_33[227]    = ( l_34 [227]);
assign l_33[228]    = ( l_34 [228]);
assign l_33[229]    = ( l_34 [229]);
assign l_33[230]    = ( l_34 [230]);
assign l_33[231]    = ( l_34 [231]);
assign l_33[232]    = ( l_34 [232]);
assign l_33[233]    = ( l_34 [233]);
assign l_33[234]    = ( l_34 [234]);
assign l_33[235]    = ( l_34 [235]);
assign l_33[236]    = ( l_34 [236]);
assign l_33[237]    = ( l_34 [237]);
assign l_33[238]    = ( l_34 [238]);
assign l_33[239]    = ( l_34 [239]);
assign l_33[240]    = ( l_34 [240]);
assign l_33[241]    = ( l_34 [241]);
assign l_33[242]    = ( l_34 [242]);
assign l_33[243]    = ( l_34 [243]);
assign l_33[244]    = ( l_34 [244]);
assign l_33[245]    = ( l_34 [245]);
assign l_33[246]    = ( l_34 [246]);
assign l_33[247]    = ( l_34 [247]);
assign l_33[248]    = ( l_34 [248]);
assign l_33[249]    = ( l_34 [249]);
assign l_33[250]    = ( l_34 [250]);
assign l_33[251]    = ( l_34 [251]);
assign l_33[252]    = ( l_34 [252]);
assign l_33[253]    = ( l_34 [253]);
assign l_33[254]    = ( l_34 [254]);
assign l_33[255]    = ( l_34 [255]);
assign l_33[256]    = ( l_34 [256]);
assign l_33[257]    = ( l_34 [257]);
assign l_33[258]    = ( l_34 [258]);
assign l_33[259]    = ( l_34 [259]);
assign l_33[260]    = ( l_34 [260]);
assign l_33[261]    = ( l_34 [261]);
assign l_33[262]    = ( l_34 [262]);
assign l_33[263]    = ( l_34 [263]);
assign l_33[264]    = ( l_34 [264]);
assign l_33[265]    = ( l_34 [265]);
assign l_33[266]    = ( l_34 [266]);
assign l_33[267]    = ( l_34 [267]);
assign l_33[268]    = ( l_34 [268]);
assign l_33[269]    = ( l_34 [269]);
assign l_33[270]    = ( l_34 [270]);
assign l_33[271]    = ( l_34 [271]);
assign l_33[272]    = ( l_34 [272]);
assign l_33[273]    = ( l_34 [273]);
assign l_33[274]    = ( l_34 [274] & !i[1818]) | ( l_34 [275] &  i[1818]);
assign l_33[275]    = ( l_34 [276] & !i[1818]) | ( l_34 [277] &  i[1818]);
assign l_33[276]    = ( l_34 [278] & !i[1818]) | ( l_34 [279] &  i[1818]);
assign l_33[277]    = ( l_34 [280] & !i[1818]) | ( l_34 [281] &  i[1818]);
assign l_33[278]    = ( l_34 [282] & !i[1818]) | ( l_34 [283] &  i[1818]);
assign l_33[279]    = ( l_34 [284] & !i[1818]) | ( l_34 [285] &  i[1818]);
assign l_33[280]    = ( l_34 [286] & !i[1818]) | ( l_34 [287] &  i[1818]);
assign l_33[281]    = ( l_34 [288] & !i[1818]) | ( l_34 [289] &  i[1818]);
assign l_33[282]    = ( l_34 [290] & !i[1818]) | ( l_34 [291] &  i[1818]);
assign l_33[283]    = ( l_34 [292] & !i[1818]) | ( l_34 [293] &  i[1818]);
assign l_33[284]    = ( l_34 [294] & !i[1818]) | ( l_34 [295] &  i[1818]);
assign l_33[285]    = ( l_34 [296] & !i[1818]) | ( l_34 [297] &  i[1818]);
assign l_33[286]    = ( l_34 [298] & !i[1818]) | ( l_34 [299] &  i[1818]);
assign l_33[287]    = ( l_34 [300] & !i[1818]) | ( l_34 [301] &  i[1818]);
assign l_33[288]    = ( l_34 [302] & !i[1818]) | ( l_34 [303] &  i[1818]);
assign l_33[289]    = ( l_34 [304] & !i[1818]) | ( l_34 [305] &  i[1818]);
assign l_33[290]    = ( l_34 [306] & !i[1818]) | ( l_34 [307] &  i[1818]);
assign l_33[291]    = ( l_34 [308] & !i[1818]) | ( l_34 [309] &  i[1818]);
assign l_33[292]    = ( l_34 [310] & !i[1818]) | ( l_34 [311] &  i[1818]);
assign l_33[293]    = ( l_34 [312] & !i[1818]) | ( l_34 [313] &  i[1818]);
assign l_33[294]    = ( l_34 [314] & !i[1818]) | ( l_34 [315] &  i[1818]);
assign l_33[295]    = ( l_34 [316] & !i[1818]) | ( l_34 [317] &  i[1818]);
assign l_33[296]    = ( l_34 [318] & !i[1818]) | ( l_34 [319] &  i[1818]);
assign l_33[297]    = ( l_34 [320] & !i[1818]) | ( l_34 [321] &  i[1818]);
assign l_33[298]    = ( l_34 [322] & !i[1818]) | ( l_34 [323] &  i[1818]);
assign l_33[299]    = ( l_34 [324] & !i[1818]) | ( l_34 [325] &  i[1818]);
assign l_33[300]    = ( l_34 [326] & !i[1818]) | ( l_34 [327] &  i[1818]);
assign l_33[301]    = ( l_34 [328] & !i[1818]) | ( l_34 [329] &  i[1818]);
assign l_33[302]    = ( l_34 [330] & !i[1818]) | ( l_34 [331] &  i[1818]);
assign l_33[303]    = ( l_34 [332] & !i[1818]) | ( l_34 [333] &  i[1818]);
assign l_33[304]    = ( l_34 [334] & !i[1818]) | ( l_34 [335] &  i[1818]);
assign l_33[305]    = ( l_34 [336] & !i[1818]) | ( l_34 [337] &  i[1818]);
assign l_33[306]    = ( l_34 [338] & !i[1818]) | ( l_34 [339] &  i[1818]);
assign l_33[307]    = ( l_34 [340] & !i[1818]) | ( l_34 [341] &  i[1818]);
assign l_33[308]    = ( l_34 [342] & !i[1818]) | ( l_34 [343] &  i[1818]);
assign l_33[309]    = ( l_34 [344] & !i[1818]) | ( l_34 [345] &  i[1818]);
assign l_33[310]    = ( l_34 [346] & !i[1818]) | ( l_34 [347] &  i[1818]);
assign l_33[311]    = ( l_34 [348] & !i[1818]) | ( l_34 [349] &  i[1818]);
assign l_33[312]    = ( l_34 [350] & !i[1818]) | ( l_34 [351] &  i[1818]);
assign l_33[313]    = ( l_34 [352] & !i[1818]) | ( l_34 [353] &  i[1818]);
assign l_33[314]    = ( l_34 [354] & !i[1818]) | ( l_34 [355] &  i[1818]);
assign l_33[315]    = ( l_34 [356] & !i[1818]) | ( l_34 [357] &  i[1818]);
assign l_33[316]    = ( l_34 [358] & !i[1818]) | ( l_34 [359] &  i[1818]);
assign l_33[317]    = ( l_34 [360] & !i[1818]) | ( l_34 [361] &  i[1818]);
assign l_33[318]    = ( l_34 [362] & !i[1818]) | ( l_34 [363] &  i[1818]);
assign l_33[319]    = ( l_34 [364] & !i[1818]) | ( l_34 [365] &  i[1818]);
assign l_33[320]    = ( l_34 [366] & !i[1818]) | ( l_34 [367] &  i[1818]);
assign l_33[321]    = ( l_34 [368] & !i[1818]) | ( l_34 [369] &  i[1818]);
assign l_33[322]    = ( l_34 [370] & !i[1818]) | ( l_34 [371] &  i[1818]);
assign l_33[323]    = ( l_34 [372] & !i[1818]) | ( l_34 [373] &  i[1818]);
assign l_33[324]    = ( l_34 [374] & !i[1818]) | ( l_34 [375] &  i[1818]);
assign l_33[325]    = ( l_34 [376] & !i[1818]) | ( l_34 [377] &  i[1818]);
assign l_33[326]    = ( l_34 [378] & !i[1818]) | ( l_34 [379] &  i[1818]);
assign l_33[327]    = ( l_34 [380] & !i[1818]) | ( l_34 [381] &  i[1818]);
assign l_33[328]    = ( l_34 [382] & !i[1818]) | ( l_34 [383] &  i[1818]);
assign l_33[329]    = ( l_34 [384] & !i[1818]) | ( l_34 [385] &  i[1818]);
assign l_33[330]    = ( l_34 [386] & !i[1818]) | ( l_34 [387] &  i[1818]);
assign l_33[331]    = ( l_34 [388] & !i[1818]) | ( l_34 [389] &  i[1818]);
assign l_33[332]    = ( l_34 [390] & !i[1818]) | ( l_34 [391] &  i[1818]);
assign l_33[333]    = ( l_34 [392] & !i[1818]) | ( l_34 [393] &  i[1818]);
assign l_33[334]    = ( l_34 [394] & !i[1818]) | ( l_34 [395] &  i[1818]);
assign l_33[335]    = ( l_34 [396] & !i[1818]) | ( l_34 [397] &  i[1818]);
assign l_33[336]    = ( l_34 [398] & !i[1818]) | ( l_34 [399] &  i[1818]);
assign l_33[337]    = ( l_34 [400] & !i[1818]) | ( l_34 [401] &  i[1818]);
assign l_33[338]    = ( l_34 [402] & !i[1818]) | ( l_34 [403] &  i[1818]);
assign l_33[339]    = ( l_34 [404] & !i[1818]) | ( l_34 [405] &  i[1818]);
assign l_33[340]    = ( l_34 [406] & !i[1818]) | ( l_34 [407] &  i[1818]);
assign l_33[341]    = ( l_34 [408] & !i[1818]) | ( l_34 [409] &  i[1818]);
assign l_33[342]    = ( l_34 [410] & !i[1818]) | ( l_34 [411] &  i[1818]);
assign l_33[343]    = ( l_34 [412] & !i[1818]) | ( l_34 [413] &  i[1818]);
assign l_33[344]    = ( l_34 [414] & !i[1818]) | ( l_34 [415] &  i[1818]);
assign l_33[345]    = ( l_34 [416] & !i[1818]) | ( l_34 [417] &  i[1818]);
assign l_33[346]    = ( l_34 [418] & !i[1818]) | ( l_34 [419] &  i[1818]);
assign l_33[347]    = ( l_34 [420] & !i[1818]) | ( l_34 [421] &  i[1818]);
assign l_33[348]    = ( l_34 [422] & !i[1818]) | ( l_34 [423] &  i[1818]);
assign l_33[349]    = ( l_34 [424] & !i[1818]) | ( l_34 [425] &  i[1818]);
assign l_33[350]    = ( l_34 [426] & !i[1818]) | ( l_34 [427] &  i[1818]);
assign l_33[351]    = ( l_34 [428] & !i[1818]) | ( l_34 [429] &  i[1818]);
assign l_33[352]    = ( l_34 [430] & !i[1818]) | ( l_34 [431] &  i[1818]);
assign l_33[353]    = ( l_34 [432] & !i[1818]) | ( l_34 [433] &  i[1818]);
assign l_33[354]    = ( l_34 [434] & !i[1818]) | ( l_34 [435] &  i[1818]);
assign l_33[355]    = ( l_34 [436] & !i[1818]) | ( l_34 [437] &  i[1818]);
assign l_33[356]    = ( l_34 [438] & !i[1818]) | ( l_34 [439] &  i[1818]);
assign l_33[357]    = ( l_34 [440] & !i[1818]) | ( l_34 [441] &  i[1818]);
assign l_33[358]    = ( l_34 [442] & !i[1818]) | ( l_34 [443] &  i[1818]);
assign l_33[359]    = ( l_34 [444] & !i[1818]) | ( l_34 [445] &  i[1818]);
assign l_33[360]    = ( l_34 [446] & !i[1818]) | ( l_34 [447] &  i[1818]);
assign l_33[361]    = ( l_34 [448] & !i[1818]) | ( l_34 [449] &  i[1818]);
assign l_33[362]    = ( l_34 [450] & !i[1818]) | ( l_34 [451] &  i[1818]);
assign l_33[363]    = ( l_34 [452] & !i[1818]) | ( l_34 [453] &  i[1818]);
assign l_33[364]    = ( l_34 [454] & !i[1818]) | ( l_34 [455] &  i[1818]);
assign l_33[365]    = ( l_34 [456] & !i[1818]) | ( l_34 [457] &  i[1818]);
assign l_33[366]    = ( l_34 [458] & !i[1818]) | ( l_34 [459] &  i[1818]);
assign l_33[367]    = ( l_34 [460] & !i[1818]) | ( l_34 [461] &  i[1818]);
assign l_33[368]    = ( l_34 [462] & !i[1818]) | ( l_34 [463] &  i[1818]);
assign l_33[369]    = ( l_34 [464] & !i[1818]) | ( l_34 [465] &  i[1818]);
assign l_33[370]    = ( l_34 [466] & !i[1818]) | ( l_34 [467] &  i[1818]);
assign l_33[371]    = ( l_34 [468] & !i[1818]) | ( l_34 [469] &  i[1818]);
assign l_33[372]    = ( l_34 [470] & !i[1818]) | ( l_34 [471] &  i[1818]);
assign l_33[373]    = ( l_34 [472] & !i[1818]) | ( l_34 [473] &  i[1818]);
assign l_33[374]    = ( l_34 [474] & !i[1818]) | ( l_34 [475] &  i[1818]);
assign l_33[375]    = ( l_34 [476] & !i[1818]) | ( l_34 [477] &  i[1818]);
assign l_33[376]    = ( l_34 [478] & !i[1818]) | ( l_34 [479] &  i[1818]);
assign l_33[377]    = ( l_34 [480] & !i[1818]) | ( l_34 [481] &  i[1818]);
assign l_33[378]    = ( l_34 [482] & !i[1818]) | ( l_34 [483] &  i[1818]);
assign l_33[379]    = ( l_34 [484] & !i[1818]) | ( l_34 [485] &  i[1818]);
assign l_33[380]    = ( l_34 [486] & !i[1818]) | ( l_34 [487] &  i[1818]);
assign l_33[381]    = ( l_34 [488] & !i[1818]) | ( l_34 [489] &  i[1818]);
assign l_33[382]    = ( l_34 [490] & !i[1818]) | ( l_34 [491] &  i[1818]);
assign l_33[383]    = ( l_34 [492] & !i[1818]) | ( l_34 [493] &  i[1818]);
assign l_33[384]    = ( l_34 [494] & !i[1818]) | ( l_34 [495] &  i[1818]);
assign l_33[385]    = ( l_34 [496] & !i[1818]) | ( l_34 [497] &  i[1818]);
assign l_33[386]    = ( l_34 [498] & !i[1818]) | ( l_34 [499] &  i[1818]);
assign l_33[387]    = ( l_34 [500] & !i[1818]) | ( l_34 [501] &  i[1818]);
assign l_33[388]    = ( l_34 [502] & !i[1818]) | ( l_34 [503] &  i[1818]);
assign l_33[389]    = ( l_34 [504] & !i[1818]) | ( l_34 [505] &  i[1818]);
assign l_33[390]    = ( l_34 [506] & !i[1818]) | ( l_34 [507] &  i[1818]);
assign l_33[391]    = ( l_34 [508] & !i[1818]) | ( l_34 [509] &  i[1818]);
assign l_33[392]    = ( l_34 [510] & !i[1818]) | ( l_34 [511] &  i[1818]);
assign l_33[393]    = ( l_34 [512] & !i[1818]) | ( l_34 [513] &  i[1818]);
assign l_33[394]    = ( l_34 [514] & !i[1818]) | ( l_34 [515] &  i[1818]);
assign l_33[395]    = ( l_34 [516] & !i[1818]) | ( l_34 [517] &  i[1818]);
assign l_33[396]    = ( l_34 [518] & !i[1818]) | ( l_34 [519] &  i[1818]);
assign l_33[397]    = ( l_34 [520] & !i[1818]) | ( l_34 [521] &  i[1818]);
assign l_33[398]    = ( l_34 [522] & !i[1818]) | ( l_34 [523] &  i[1818]);
assign l_33[399]    = ( l_34 [524] & !i[1818]) | ( l_34 [525] &  i[1818]);
assign l_33[400]    = ( l_34 [526] & !i[1818]) | ( l_34 [527] &  i[1818]);
assign l_33[401]    = ( l_34 [528] & !i[1818]) | ( l_34 [529] &  i[1818]);
assign l_34[0]    = ( l_35 [0]);
assign l_34[1]    = ( l_35 [1] & !i[1813]);
assign l_34[2]    = ( l_35 [2] & !i[1813]);
assign l_34[3]    = (!i[1813]) | ( l_35 [3] &  i[1813]);
assign l_34[4]    = (!i[1813]) | ( l_35 [4] &  i[1813]);
assign l_34[5]    = ( l_35 [5] & !i[1813]);
assign l_34[6]    = ( l_35 [6] & !i[1813]);
assign l_34[7]    = (!i[1813]) | ( l_35 [7] &  i[1813]);
assign l_34[8]    = (!i[1813]) | ( l_35 [8] &  i[1813]);
assign l_34[9]    = ( l_35 [9] & !i[1813]) | ( l_35 [10] &  i[1813]);
assign l_34[10]    = ( l_35 [10]);
assign l_34[11]    = ( l_35 [11] & !i[1813]) | ( l_35 [10] &  i[1813]);
assign l_34[12]    = ( l_35 [10] & !i[1813]) | ( l_35 [12] &  i[1813]);
assign l_34[13]    = ( l_35 [10] & !i[1813]) | ( l_35 [13] &  i[1813]);
assign l_34[14]    = ( l_35 [14] & !i[1813]) | ( l_35 [10] &  i[1813]);
assign l_34[15]    = ( l_35 [15] & !i[1813]) | ( l_35 [10] &  i[1813]);
assign l_34[16]    = ( l_35 [10] & !i[1813]) | ( l_35 [16] &  i[1813]);
assign l_34[17]    = ( l_35 [10] & !i[1813]) | ( l_35 [17] &  i[1813]);
assign l_34[18]    = ( l_35 [18] & !i[1813]) | ( l_35 [19] &  i[1813]);
assign l_34[19]    = ( l_35 [20] & !i[1813]) | ( l_35 [21] &  i[1813]);
assign l_34[20]    = ( l_35 [22] & !i[1813]) | ( l_35 [23] &  i[1813]);
assign l_34[21]    = ( l_35 [24] & !i[1813]) | ( l_35 [25] &  i[1813]);
assign l_34[22]    = ( l_35 [26] & !i[1813]) | ( l_35 [27] &  i[1813]);
assign l_34[23]    = ( l_35 [28] & !i[1813]) | ( l_35 [29] &  i[1813]);
assign l_34[24]    = ( l_35 [30] & !i[1813]) | ( l_35 [31] &  i[1813]);
assign l_34[25]    = ( l_35 [32] & !i[1813]) | ( l_35 [33] &  i[1813]);
assign l_34[26]    = ( l_35 [34] & !i[1813]) | ( l_35 [35] &  i[1813]);
assign l_34[27]    = ( l_35 [36] & !i[1813]) | ( l_35 [37] &  i[1813]);
assign l_34[28]    = ( l_35 [38] & !i[1813]) | ( l_35 [39] &  i[1813]);
assign l_34[29]    = ( l_35 [40] & !i[1813]) | ( l_35 [41] &  i[1813]);
assign l_34[30]    = ( l_35 [42] & !i[1813]) | ( l_35 [43] &  i[1813]);
assign l_34[31]    = ( l_35 [44] & !i[1813]) | ( l_35 [45] &  i[1813]);
assign l_34[32]    = ( l_35 [46] & !i[1813]) | ( l_35 [47] &  i[1813]);
assign l_34[33]    = ( l_35 [48] & !i[1813]) | ( l_35 [49] &  i[1813]);
assign l_34[34]    = ( l_35 [50] & !i[1813]) | ( l_35 [51] &  i[1813]);
assign l_34[35]    = ( l_35 [52] & !i[1813]) | ( l_35 [53] &  i[1813]);
assign l_34[36]    = ( l_35 [54] & !i[1813]) | ( l_35 [55] &  i[1813]);
assign l_34[37]    = ( l_35 [56] & !i[1813]) | ( l_35 [57] &  i[1813]);
assign l_34[38]    = ( l_35 [58] & !i[1813]) | ( l_35 [59] &  i[1813]);
assign l_34[39]    = ( l_35 [60] & !i[1813]) | ( l_35 [61] &  i[1813]);
assign l_34[40]    = ( l_35 [62] & !i[1813]) | ( l_35 [63] &  i[1813]);
assign l_34[41]    = ( l_35 [64] & !i[1813]) | ( l_35 [65] &  i[1813]);
assign l_34[42]    = ( l_35 [66] & !i[1813]) | ( l_35 [67] &  i[1813]);
assign l_34[43]    = ( l_35 [68] & !i[1813]) | ( l_35 [69] &  i[1813]);
assign l_34[44]    = ( l_35 [70] & !i[1813]) | ( l_35 [71] &  i[1813]);
assign l_34[45]    = ( l_35 [72] & !i[1813]) | ( l_35 [73] &  i[1813]);
assign l_34[46]    = ( l_35 [74] & !i[1813]) | ( l_35 [75] &  i[1813]);
assign l_34[47]    = ( l_35 [76] & !i[1813]) | ( l_35 [77] &  i[1813]);
assign l_34[48]    = ( l_35 [78] & !i[1813]) | ( l_35 [79] &  i[1813]);
assign l_34[49]    = ( l_35 [80] & !i[1813]) | ( l_35 [81] &  i[1813]);
assign l_34[50]    = ( l_35 [82] & !i[1813]) | ( l_35 [83] &  i[1813]);
assign l_34[51]    = ( l_35 [84] & !i[1813]) | ( l_35 [85] &  i[1813]);
assign l_34[52]    = ( l_35 [86] & !i[1813]) | ( l_35 [87] &  i[1813]);
assign l_34[53]    = ( l_35 [88] & !i[1813]) | ( l_35 [89] &  i[1813]);
assign l_34[54]    = ( l_35 [90] & !i[1813]) | ( l_35 [91] &  i[1813]);
assign l_34[55]    = ( l_35 [92] & !i[1813]) | ( l_35 [93] &  i[1813]);
assign l_34[56]    = ( l_35 [94] & !i[1813]) | ( l_35 [95] &  i[1813]);
assign l_34[57]    = ( l_35 [96] & !i[1813]) | ( l_35 [97] &  i[1813]);
assign l_34[58]    = ( l_35 [98] & !i[1813]) | ( l_35 [99] &  i[1813]);
assign l_34[59]    = ( l_35 [100] & !i[1813]) | ( l_35 [101] &  i[1813]);
assign l_34[60]    = ( l_35 [102] & !i[1813]) | ( l_35 [103] &  i[1813]);
assign l_34[61]    = ( l_35 [104] & !i[1813]) | ( l_35 [105] &  i[1813]);
assign l_34[62]    = ( l_35 [106] & !i[1813]) | ( l_35 [107] &  i[1813]);
assign l_34[63]    = ( l_35 [108] & !i[1813]) | ( l_35 [109] &  i[1813]);
assign l_34[64]    = ( l_35 [110] & !i[1813]) | ( l_35 [111] &  i[1813]);
assign l_34[65]    = ( l_35 [112] & !i[1813]) | ( l_35 [113] &  i[1813]);
assign l_34[66]    = ( l_35 [114] & !i[1813]) | ( l_35 [115] &  i[1813]);
assign l_34[67]    = ( l_35 [116] & !i[1813]) | ( l_35 [117] &  i[1813]);
assign l_34[68]    = ( l_35 [118] & !i[1813]) | ( l_35 [119] &  i[1813]);
assign l_34[69]    = ( l_35 [120] & !i[1813]) | ( l_35 [121] &  i[1813]);
assign l_34[70]    = ( l_35 [122] & !i[1813]) | ( l_35 [123] &  i[1813]);
assign l_34[71]    = ( l_35 [124] & !i[1813]) | ( l_35 [125] &  i[1813]);
assign l_34[72]    = ( l_35 [126] & !i[1813]) | ( l_35 [127] &  i[1813]);
assign l_34[73]    = ( l_35 [128] & !i[1813]) | ( l_35 [129] &  i[1813]);
assign l_34[74]    = ( l_35 [130] & !i[1813]) | ( l_35 [131] &  i[1813]);
assign l_34[75]    = ( l_35 [132] & !i[1813]) | ( l_35 [133] &  i[1813]);
assign l_34[76]    = ( l_35 [134] & !i[1813]) | ( l_35 [135] &  i[1813]);
assign l_34[77]    = ( l_35 [136] & !i[1813]) | ( l_35 [137] &  i[1813]);
assign l_34[78]    = ( l_35 [138] & !i[1813]) | ( l_35 [139] &  i[1813]);
assign l_34[79]    = ( l_35 [140] & !i[1813]) | ( l_35 [141] &  i[1813]);
assign l_34[80]    = ( l_35 [142] & !i[1813]) | ( l_35 [143] &  i[1813]);
assign l_34[81]    = ( l_35 [144] & !i[1813]) | ( l_35 [145] &  i[1813]);
assign l_34[82]    = ( l_35 [146] & !i[1813]) | ( l_35 [147] &  i[1813]);
assign l_34[83]    = ( l_35 [148] & !i[1813]) | ( l_35 [149] &  i[1813]);
assign l_34[84]    = ( l_35 [150] & !i[1813]) | ( l_35 [151] &  i[1813]);
assign l_34[85]    = ( l_35 [152] & !i[1813]) | ( l_35 [153] &  i[1813]);
assign l_34[86]    = ( l_35 [154] & !i[1813]) | ( l_35 [155] &  i[1813]);
assign l_34[87]    = ( l_35 [156] & !i[1813]) | ( l_35 [157] &  i[1813]);
assign l_34[88]    = ( l_35 [158] & !i[1813]) | ( l_35 [159] &  i[1813]);
assign l_34[89]    = ( l_35 [160] & !i[1813]) | ( l_35 [161] &  i[1813]);
assign l_34[90]    = ( l_35 [162] & !i[1813]) | ( l_35 [163] &  i[1813]);
assign l_34[91]    = ( l_35 [164] & !i[1813]) | ( l_35 [165] &  i[1813]);
assign l_34[92]    = ( l_35 [166] & !i[1813]) | ( l_35 [167] &  i[1813]);
assign l_34[93]    = ( l_35 [168] & !i[1813]) | ( l_35 [169] &  i[1813]);
assign l_34[94]    = ( l_35 [170] & !i[1813]) | ( l_35 [171] &  i[1813]);
assign l_34[95]    = ( l_35 [172] & !i[1813]) | ( l_35 [173] &  i[1813]);
assign l_34[96]    = ( l_35 [174] & !i[1813]) | ( l_35 [175] &  i[1813]);
assign l_34[97]    = ( l_35 [176] & !i[1813]) | ( l_35 [177] &  i[1813]);
assign l_34[98]    = ( l_35 [178] & !i[1813]) | ( l_35 [179] &  i[1813]);
assign l_34[99]    = ( l_35 [180] & !i[1813]) | ( l_35 [181] &  i[1813]);
assign l_34[100]    = ( l_35 [182] & !i[1813]) | ( l_35 [183] &  i[1813]);
assign l_34[101]    = ( l_35 [184] & !i[1813]) | ( l_35 [185] &  i[1813]);
assign l_34[102]    = ( l_35 [186] & !i[1813]) | ( l_35 [187] &  i[1813]);
assign l_34[103]    = ( l_35 [188] & !i[1813]) | ( l_35 [189] &  i[1813]);
assign l_34[104]    = ( l_35 [190] & !i[1813]) | ( l_35 [191] &  i[1813]);
assign l_34[105]    = ( l_35 [192] & !i[1813]) | ( l_35 [193] &  i[1813]);
assign l_34[106]    = ( l_35 [194] & !i[1813]) | ( l_35 [195] &  i[1813]);
assign l_34[107]    = ( l_35 [196] & !i[1813]) | ( l_35 [197] &  i[1813]);
assign l_34[108]    = ( l_35 [198] & !i[1813]) | ( l_35 [199] &  i[1813]);
assign l_34[109]    = ( l_35 [200] & !i[1813]) | ( l_35 [201] &  i[1813]);
assign l_34[110]    = ( l_35 [202] & !i[1813]) | ( l_35 [203] &  i[1813]);
assign l_34[111]    = ( l_35 [204] & !i[1813]) | ( l_35 [205] &  i[1813]);
assign l_34[112]    = ( l_35 [206] & !i[1813]) | ( l_35 [207] &  i[1813]);
assign l_34[113]    = ( l_35 [208] & !i[1813]) | ( l_35 [209] &  i[1813]);
assign l_34[114]    = ( l_35 [210] & !i[1813]) | ( l_35 [211] &  i[1813]);
assign l_34[115]    = ( l_35 [212] & !i[1813]) | ( l_35 [213] &  i[1813]);
assign l_34[116]    = ( l_35 [214] & !i[1813]) | ( l_35 [215] &  i[1813]);
assign l_34[117]    = ( l_35 [216] & !i[1813]) | ( l_35 [217] &  i[1813]);
assign l_34[118]    = ( l_35 [218] & !i[1813]) | ( l_35 [219] &  i[1813]);
assign l_34[119]    = ( l_35 [220] & !i[1813]) | ( l_35 [221] &  i[1813]);
assign l_34[120]    = ( l_35 [222] & !i[1813]) | ( l_35 [223] &  i[1813]);
assign l_34[121]    = ( l_35 [224] & !i[1813]) | ( l_35 [225] &  i[1813]);
assign l_34[122]    = ( l_35 [226] & !i[1813]) | ( l_35 [227] &  i[1813]);
assign l_34[123]    = ( l_35 [228] & !i[1813]) | ( l_35 [229] &  i[1813]);
assign l_34[124]    = ( l_35 [230] & !i[1813]) | ( l_35 [231] &  i[1813]);
assign l_34[125]    = ( l_35 [232] & !i[1813]) | ( l_35 [233] &  i[1813]);
assign l_34[126]    = ( l_35 [234] & !i[1813]) | ( l_35 [235] &  i[1813]);
assign l_34[127]    = ( l_35 [236] & !i[1813]) | ( l_35 [237] &  i[1813]);
assign l_34[128]    = ( l_35 [238] & !i[1813]) | ( l_35 [239] &  i[1813]);
assign l_34[129]    = ( l_35 [240] & !i[1813]) | ( l_35 [241] &  i[1813]);
assign l_34[130]    = ( l_35 [242] & !i[1813]) | ( l_35 [243] &  i[1813]);
assign l_34[131]    = ( l_35 [244] & !i[1813]) | ( l_35 [245] &  i[1813]);
assign l_34[132]    = ( l_35 [246] & !i[1813]) | ( l_35 [247] &  i[1813]);
assign l_34[133]    = ( l_35 [248] & !i[1813]) | ( l_35 [249] &  i[1813]);
assign l_34[134]    = ( l_35 [250] & !i[1813]) | ( l_35 [251] &  i[1813]);
assign l_34[135]    = ( l_35 [252] & !i[1813]) | ( l_35 [253] &  i[1813]);
assign l_34[136]    = ( l_35 [254] & !i[1813]) | ( l_35 [255] &  i[1813]);
assign l_34[137]    = ( l_35 [256] & !i[1813]) | ( l_35 [257] &  i[1813]);
assign l_34[138]    = ( l_35 [258] & !i[1813]) | ( l_35 [259] &  i[1813]);
assign l_34[139]    = ( l_35 [260] & !i[1813]) | ( l_35 [261] &  i[1813]);
assign l_34[140]    = ( l_35 [262] & !i[1813]) | ( l_35 [263] &  i[1813]);
assign l_34[141]    = ( l_35 [264] & !i[1813]) | ( l_35 [265] &  i[1813]);
assign l_34[142]    = ( l_35 [266] & !i[1813]) | ( l_35 [267] &  i[1813]);
assign l_34[143]    = ( l_35 [268] & !i[1813]) | ( l_35 [269] &  i[1813]);
assign l_34[144]    = ( l_35 [270] & !i[1813]) | ( l_35 [271] &  i[1813]);
assign l_34[145]    = ( l_35 [272] & !i[1813]) | ( l_35 [273] &  i[1813]);
assign l_34[146]    = ( l_35 [274] & !i[1813]) | ( l_35 [275] &  i[1813]);
assign l_34[147]    = ( l_35 [276] & !i[1813]) | ( l_35 [277] &  i[1813]);
assign l_34[148]    = ( l_35 [278] & !i[1813]) | ( l_35 [279] &  i[1813]);
assign l_34[149]    = ( l_35 [280] & !i[1813]) | ( l_35 [281] &  i[1813]);
assign l_34[150]    = ( l_35 [282] & !i[1813]) | ( l_35 [283] &  i[1813]);
assign l_34[151]    = ( l_35 [284] & !i[1813]) | ( l_35 [285] &  i[1813]);
assign l_34[152]    = ( l_35 [286] & !i[1813]) | ( l_35 [287] &  i[1813]);
assign l_34[153]    = ( l_35 [288] & !i[1813]) | ( l_35 [289] &  i[1813]);
assign l_34[154]    = ( l_35 [290] & !i[1813]) | ( l_35 [291] &  i[1813]);
assign l_34[155]    = ( l_35 [292] & !i[1813]) | ( l_35 [293] &  i[1813]);
assign l_34[156]    = ( l_35 [294] & !i[1813]) | ( l_35 [295] &  i[1813]);
assign l_34[157]    = ( l_35 [296] & !i[1813]) | ( l_35 [297] &  i[1813]);
assign l_34[158]    = ( l_35 [298] & !i[1813]) | ( l_35 [299] &  i[1813]);
assign l_34[159]    = ( l_35 [300] & !i[1813]) | ( l_35 [301] &  i[1813]);
assign l_34[160]    = ( l_35 [302] & !i[1813]) | ( l_35 [303] &  i[1813]);
assign l_34[161]    = ( l_35 [304] & !i[1813]) | ( l_35 [305] &  i[1813]);
assign l_34[162]    = ( l_35 [306] & !i[1813]) | ( l_35 [307] &  i[1813]);
assign l_34[163]    = ( l_35 [308] & !i[1813]) | ( l_35 [309] &  i[1813]);
assign l_34[164]    = ( l_35 [310] & !i[1813]) | ( l_35 [311] &  i[1813]);
assign l_34[165]    = ( l_35 [312] & !i[1813]) | ( l_35 [313] &  i[1813]);
assign l_34[166]    = ( l_35 [314] & !i[1813]) | ( l_35 [315] &  i[1813]);
assign l_34[167]    = ( l_35 [316] & !i[1813]) | ( l_35 [317] &  i[1813]);
assign l_34[168]    = ( l_35 [318] & !i[1813]) | ( l_35 [319] &  i[1813]);
assign l_34[169]    = ( l_35 [320] & !i[1813]) | ( l_35 [321] &  i[1813]);
assign l_34[170]    = ( l_35 [322] & !i[1813]) | ( l_35 [323] &  i[1813]);
assign l_34[171]    = ( l_35 [324] & !i[1813]) | ( l_35 [325] &  i[1813]);
assign l_34[172]    = ( l_35 [326] & !i[1813]) | ( l_35 [327] &  i[1813]);
assign l_34[173]    = ( l_35 [328] & !i[1813]) | ( l_35 [329] &  i[1813]);
assign l_34[174]    = ( l_35 [330] & !i[1813]) | ( l_35 [331] &  i[1813]);
assign l_34[175]    = ( l_35 [332] & !i[1813]) | ( l_35 [333] &  i[1813]);
assign l_34[176]    = ( l_35 [334] & !i[1813]) | ( l_35 [335] &  i[1813]);
assign l_34[177]    = ( l_35 [336] & !i[1813]) | ( l_35 [337] &  i[1813]);
assign l_34[178]    = ( l_35 [338] & !i[1813]) | ( l_35 [339] &  i[1813]);
assign l_34[179]    = ( l_35 [340] & !i[1813]) | ( l_35 [341] &  i[1813]);
assign l_34[180]    = ( l_35 [342] & !i[1813]) | ( l_35 [343] &  i[1813]);
assign l_34[181]    = ( l_35 [344] & !i[1813]) | ( l_35 [345] &  i[1813]);
assign l_34[182]    = ( l_35 [346] & !i[1813]) | ( l_35 [347] &  i[1813]);
assign l_34[183]    = ( l_35 [348] & !i[1813]) | ( l_35 [349] &  i[1813]);
assign l_34[184]    = ( l_35 [350] & !i[1813]) | ( l_35 [351] &  i[1813]);
assign l_34[185]    = ( l_35 [352] & !i[1813]) | ( l_35 [353] &  i[1813]);
assign l_34[186]    = ( l_35 [354] & !i[1813]) | ( l_35 [355] &  i[1813]);
assign l_34[187]    = ( l_35 [356] & !i[1813]) | ( l_35 [357] &  i[1813]);
assign l_34[188]    = ( l_35 [358] & !i[1813]) | ( l_35 [359] &  i[1813]);
assign l_34[189]    = ( l_35 [360] & !i[1813]) | ( l_35 [361] &  i[1813]);
assign l_34[190]    = ( l_35 [362] & !i[1813]) | ( l_35 [363] &  i[1813]);
assign l_34[191]    = ( l_35 [364] & !i[1813]) | ( l_35 [365] &  i[1813]);
assign l_34[192]    = ( l_35 [366] & !i[1813]) | ( l_35 [367] &  i[1813]);
assign l_34[193]    = ( l_35 [368] & !i[1813]) | ( l_35 [369] &  i[1813]);
assign l_34[194]    = ( l_35 [370] & !i[1813]) | ( l_35 [371] &  i[1813]);
assign l_34[195]    = ( l_35 [372] & !i[1813]) | ( l_35 [373] &  i[1813]);
assign l_34[196]    = ( l_35 [374] & !i[1813]) | ( l_35 [375] &  i[1813]);
assign l_34[197]    = ( l_35 [376] & !i[1813]) | ( l_35 [377] &  i[1813]);
assign l_34[198]    = ( l_35 [378] & !i[1813]) | ( l_35 [379] &  i[1813]);
assign l_34[199]    = ( l_35 [380] & !i[1813]) | ( l_35 [381] &  i[1813]);
assign l_34[200]    = ( l_35 [382] & !i[1813]) | ( l_35 [383] &  i[1813]);
assign l_34[201]    = ( l_35 [384] & !i[1813]) | ( l_35 [385] &  i[1813]);
assign l_34[202]    = ( l_35 [386] & !i[1813]) | ( l_35 [387] &  i[1813]);
assign l_34[203]    = ( l_35 [388] & !i[1813]) | ( l_35 [389] &  i[1813]);
assign l_34[204]    = ( l_35 [390] & !i[1813]) | ( l_35 [391] &  i[1813]);
assign l_34[205]    = ( l_35 [392] & !i[1813]) | ( l_35 [393] &  i[1813]);
assign l_34[206]    = ( l_35 [394] & !i[1813]) | ( l_35 [395] &  i[1813]);
assign l_34[207]    = ( l_35 [396] & !i[1813]) | ( l_35 [397] &  i[1813]);
assign l_34[208]    = ( l_35 [398] & !i[1813]) | ( l_35 [399] &  i[1813]);
assign l_34[209]    = ( l_35 [400] & !i[1813]) | ( l_35 [401] &  i[1813]);
assign l_34[210]    = ( l_35 [402] & !i[1813]) | ( l_35 [403] &  i[1813]);
assign l_34[211]    = ( l_35 [404] & !i[1813]) | ( l_35 [405] &  i[1813]);
assign l_34[212]    = ( l_35 [406] & !i[1813]) | ( l_35 [407] &  i[1813]);
assign l_34[213]    = ( l_35 [408] & !i[1813]) | ( l_35 [409] &  i[1813]);
assign l_34[214]    = ( l_35 [410] & !i[1813]) | ( l_35 [411] &  i[1813]);
assign l_34[215]    = ( l_35 [412] & !i[1813]) | ( l_35 [413] &  i[1813]);
assign l_34[216]    = ( l_35 [414] & !i[1813]) | ( l_35 [415] &  i[1813]);
assign l_34[217]    = ( l_35 [416] & !i[1813]) | ( l_35 [417] &  i[1813]);
assign l_34[218]    = ( l_35 [418] & !i[1813]) | ( l_35 [419] &  i[1813]);
assign l_34[219]    = ( l_35 [420] & !i[1813]) | ( l_35 [421] &  i[1813]);
assign l_34[220]    = ( l_35 [422] & !i[1813]) | ( l_35 [423] &  i[1813]);
assign l_34[221]    = ( l_35 [424] & !i[1813]) | ( l_35 [425] &  i[1813]);
assign l_34[222]    = ( l_35 [426] & !i[1813]) | ( l_35 [427] &  i[1813]);
assign l_34[223]    = ( l_35 [428] & !i[1813]) | ( l_35 [429] &  i[1813]);
assign l_34[224]    = ( l_35 [430] & !i[1813]) | ( l_35 [431] &  i[1813]);
assign l_34[225]    = ( l_35 [432] & !i[1813]) | ( l_35 [433] &  i[1813]);
assign l_34[226]    = ( l_35 [434] & !i[1813]) | ( l_35 [435] &  i[1813]);
assign l_34[227]    = ( l_35 [436] & !i[1813]) | ( l_35 [437] &  i[1813]);
assign l_34[228]    = ( l_35 [438] & !i[1813]) | ( l_35 [439] &  i[1813]);
assign l_34[229]    = ( l_35 [440] & !i[1813]) | ( l_35 [441] &  i[1813]);
assign l_34[230]    = ( l_35 [442] & !i[1813]) | ( l_35 [443] &  i[1813]);
assign l_34[231]    = ( l_35 [444] & !i[1813]) | ( l_35 [445] &  i[1813]);
assign l_34[232]    = ( l_35 [446] & !i[1813]) | ( l_35 [447] &  i[1813]);
assign l_34[233]    = ( l_35 [448] & !i[1813]) | ( l_35 [449] &  i[1813]);
assign l_34[234]    = ( l_35 [450] & !i[1813]) | ( l_35 [451] &  i[1813]);
assign l_34[235]    = ( l_35 [452] & !i[1813]) | ( l_35 [453] &  i[1813]);
assign l_34[236]    = ( l_35 [454] & !i[1813]) | ( l_35 [455] &  i[1813]);
assign l_34[237]    = ( l_35 [456] & !i[1813]) | ( l_35 [457] &  i[1813]);
assign l_34[238]    = ( l_35 [458] & !i[1813]) | ( l_35 [459] &  i[1813]);
assign l_34[239]    = ( l_35 [460] & !i[1813]) | ( l_35 [461] &  i[1813]);
assign l_34[240]    = ( l_35 [462] & !i[1813]) | ( l_35 [463] &  i[1813]);
assign l_34[241]    = ( l_35 [464] & !i[1813]) | ( l_35 [465] &  i[1813]);
assign l_34[242]    = ( l_35 [466] & !i[1813]) | ( l_35 [467] &  i[1813]);
assign l_34[243]    = ( l_35 [468] & !i[1813]) | ( l_35 [469] &  i[1813]);
assign l_34[244]    = ( l_35 [470] & !i[1813]) | ( l_35 [471] &  i[1813]);
assign l_34[245]    = ( l_35 [472] & !i[1813]) | ( l_35 [473] &  i[1813]);
assign l_34[246]    = ( l_35 [474] & !i[1813]) | ( l_35 [475] &  i[1813]);
assign l_34[247]    = ( l_35 [476] & !i[1813]) | ( l_35 [477] &  i[1813]);
assign l_34[248]    = ( l_35 [478] & !i[1813]) | ( l_35 [479] &  i[1813]);
assign l_34[249]    = ( l_35 [480] & !i[1813]) | ( l_35 [481] &  i[1813]);
assign l_34[250]    = ( l_35 [482] & !i[1813]) | ( l_35 [483] &  i[1813]);
assign l_34[251]    = ( l_35 [484] & !i[1813]) | ( l_35 [485] &  i[1813]);
assign l_34[252]    = ( l_35 [486] & !i[1813]) | ( l_35 [487] &  i[1813]);
assign l_34[253]    = ( l_35 [488] & !i[1813]) | ( l_35 [489] &  i[1813]);
assign l_34[254]    = ( l_35 [490] & !i[1813]) | ( l_35 [491] &  i[1813]);
assign l_34[255]    = ( l_35 [492] & !i[1813]) | ( l_35 [493] &  i[1813]);
assign l_34[256]    = ( l_35 [494] & !i[1813]) | ( l_35 [495] &  i[1813]);
assign l_34[257]    = ( l_35 [496] & !i[1813]) | ( l_35 [497] &  i[1813]);
assign l_34[258]    = ( l_35 [498] & !i[1813]) | ( l_35 [499] &  i[1813]);
assign l_34[259]    = ( l_35 [500] & !i[1813]) | ( l_35 [501] &  i[1813]);
assign l_34[260]    = ( l_35 [502] & !i[1813]) | ( l_35 [503] &  i[1813]);
assign l_34[261]    = ( l_35 [504] & !i[1813]) | ( l_35 [505] &  i[1813]);
assign l_34[262]    = ( l_35 [506] & !i[1813]) | ( l_35 [507] &  i[1813]);
assign l_34[263]    = ( l_35 [508] & !i[1813]) | ( l_35 [509] &  i[1813]);
assign l_34[264]    = ( l_35 [510] & !i[1813]) | ( l_35 [511] &  i[1813]);
assign l_34[265]    = ( l_35 [512] & !i[1813]) | ( l_35 [513] &  i[1813]);
assign l_34[266]    = ( l_35 [514] & !i[1813]) | ( l_35 [515] &  i[1813]);
assign l_34[267]    = ( l_35 [516] & !i[1813]) | ( l_35 [517] &  i[1813]);
assign l_34[268]    = ( l_35 [518] & !i[1813]) | ( l_35 [519] &  i[1813]);
assign l_34[269]    = ( l_35 [520] & !i[1813]) | ( l_35 [521] &  i[1813]);
assign l_34[270]    = ( l_35 [522] & !i[1813]) | ( l_35 [523] &  i[1813]);
assign l_34[271]    = ( l_35 [524] & !i[1813]) | ( l_35 [525] &  i[1813]);
assign l_34[272]    = ( l_35 [526] & !i[1813]) | ( l_35 [527] &  i[1813]);
assign l_34[273]    = ( l_35 [528] & !i[1813]) | ( l_35 [529] &  i[1813]);
assign l_34[274]    = ( l_35 [530]);
assign l_34[275]    = ( l_35 [531]);
assign l_34[276]    = ( l_35 [532]);
assign l_34[277]    = ( l_35 [533]);
assign l_34[278]    = ( l_35 [534]);
assign l_34[279]    = ( l_35 [535]);
assign l_34[280]    = ( l_35 [536]);
assign l_34[281]    = ( l_35 [537]);
assign l_34[282]    = ( l_35 [538]);
assign l_34[283]    = ( l_35 [539]);
assign l_34[284]    = ( l_35 [540]);
assign l_34[285]    = ( l_35 [541]);
assign l_34[286]    = ( l_35 [542]);
assign l_34[287]    = ( l_35 [543]);
assign l_34[288]    = ( l_35 [544]);
assign l_34[289]    = ( l_35 [545]);
assign l_34[290]    = ( l_35 [546]);
assign l_34[291]    = ( l_35 [547]);
assign l_34[292]    = ( l_35 [548]);
assign l_34[293]    = ( l_35 [549]);
assign l_34[294]    = ( l_35 [550]);
assign l_34[295]    = ( l_35 [551]);
assign l_34[296]    = ( l_35 [552]);
assign l_34[297]    = ( l_35 [553]);
assign l_34[298]    = ( l_35 [554]);
assign l_34[299]    = ( l_35 [555]);
assign l_34[300]    = ( l_35 [556]);
assign l_34[301]    = ( l_35 [557]);
assign l_34[302]    = ( l_35 [558]);
assign l_34[303]    = ( l_35 [559]);
assign l_34[304]    = ( l_35 [560]);
assign l_34[305]    = ( l_35 [561]);
assign l_34[306]    = ( l_35 [562]);
assign l_34[307]    = ( l_35 [563]);
assign l_34[308]    = ( l_35 [564]);
assign l_34[309]    = ( l_35 [565]);
assign l_34[310]    = ( l_35 [566]);
assign l_34[311]    = ( l_35 [567]);
assign l_34[312]    = ( l_35 [568]);
assign l_34[313]    = ( l_35 [569]);
assign l_34[314]    = ( l_35 [570]);
assign l_34[315]    = ( l_35 [571]);
assign l_34[316]    = ( l_35 [572]);
assign l_34[317]    = ( l_35 [573]);
assign l_34[318]    = ( l_35 [574]);
assign l_34[319]    = ( l_35 [575]);
assign l_34[320]    = ( l_35 [576]);
assign l_34[321]    = ( l_35 [577]);
assign l_34[322]    = ( l_35 [578]);
assign l_34[323]    = ( l_35 [579]);
assign l_34[324]    = ( l_35 [580]);
assign l_34[325]    = ( l_35 [581]);
assign l_34[326]    = ( l_35 [582]);
assign l_34[327]    = ( l_35 [583]);
assign l_34[328]    = ( l_35 [584]);
assign l_34[329]    = ( l_35 [585]);
assign l_34[330]    = ( l_35 [586]);
assign l_34[331]    = ( l_35 [587]);
assign l_34[332]    = ( l_35 [588]);
assign l_34[333]    = ( l_35 [589]);
assign l_34[334]    = ( l_35 [590]);
assign l_34[335]    = ( l_35 [591]);
assign l_34[336]    = ( l_35 [592]);
assign l_34[337]    = ( l_35 [593]);
assign l_34[338]    = ( l_35 [594]);
assign l_34[339]    = ( l_35 [595]);
assign l_34[340]    = ( l_35 [596]);
assign l_34[341]    = ( l_35 [597]);
assign l_34[342]    = ( l_35 [598]);
assign l_34[343]    = ( l_35 [599]);
assign l_34[344]    = ( l_35 [600]);
assign l_34[345]    = ( l_35 [601]);
assign l_34[346]    = ( l_35 [602]);
assign l_34[347]    = ( l_35 [603]);
assign l_34[348]    = ( l_35 [604]);
assign l_34[349]    = ( l_35 [605]);
assign l_34[350]    = ( l_35 [606]);
assign l_34[351]    = ( l_35 [607]);
assign l_34[352]    = ( l_35 [608]);
assign l_34[353]    = ( l_35 [609]);
assign l_34[354]    = ( l_35 [610]);
assign l_34[355]    = ( l_35 [611]);
assign l_34[356]    = ( l_35 [612]);
assign l_34[357]    = ( l_35 [613]);
assign l_34[358]    = ( l_35 [614]);
assign l_34[359]    = ( l_35 [615]);
assign l_34[360]    = ( l_35 [616]);
assign l_34[361]    = ( l_35 [617]);
assign l_34[362]    = ( l_35 [618]);
assign l_34[363]    = ( l_35 [619]);
assign l_34[364]    = ( l_35 [620]);
assign l_34[365]    = ( l_35 [621]);
assign l_34[366]    = ( l_35 [622]);
assign l_34[367]    = ( l_35 [623]);
assign l_34[368]    = ( l_35 [624]);
assign l_34[369]    = ( l_35 [625]);
assign l_34[370]    = ( l_35 [626]);
assign l_34[371]    = ( l_35 [627]);
assign l_34[372]    = ( l_35 [628]);
assign l_34[373]    = ( l_35 [629]);
assign l_34[374]    = ( l_35 [630]);
assign l_34[375]    = ( l_35 [631]);
assign l_34[376]    = ( l_35 [632]);
assign l_34[377]    = ( l_35 [633]);
assign l_34[378]    = ( l_35 [634]);
assign l_34[379]    = ( l_35 [635]);
assign l_34[380]    = ( l_35 [636]);
assign l_34[381]    = ( l_35 [637]);
assign l_34[382]    = ( l_35 [638]);
assign l_34[383]    = ( l_35 [639]);
assign l_34[384]    = ( l_35 [640]);
assign l_34[385]    = ( l_35 [641]);
assign l_34[386]    = ( l_35 [642]);
assign l_34[387]    = ( l_35 [643]);
assign l_34[388]    = ( l_35 [644]);
assign l_34[389]    = ( l_35 [645]);
assign l_34[390]    = ( l_35 [646]);
assign l_34[391]    = ( l_35 [647]);
assign l_34[392]    = ( l_35 [648]);
assign l_34[393]    = ( l_35 [649]);
assign l_34[394]    = ( l_35 [650]);
assign l_34[395]    = ( l_35 [651]);
assign l_34[396]    = ( l_35 [652]);
assign l_34[397]    = ( l_35 [653]);
assign l_34[398]    = ( l_35 [654]);
assign l_34[399]    = ( l_35 [655]);
assign l_34[400]    = ( l_35 [656]);
assign l_34[401]    = ( l_35 [657]);
assign l_34[402]    = ( l_35 [658]);
assign l_34[403]    = ( l_35 [659]);
assign l_34[404]    = ( l_35 [660]);
assign l_34[405]    = ( l_35 [661]);
assign l_34[406]    = ( l_35 [662]);
assign l_34[407]    = ( l_35 [663]);
assign l_34[408]    = ( l_35 [664]);
assign l_34[409]    = ( l_35 [665]);
assign l_34[410]    = ( l_35 [666]);
assign l_34[411]    = ( l_35 [667]);
assign l_34[412]    = ( l_35 [668]);
assign l_34[413]    = ( l_35 [669]);
assign l_34[414]    = ( l_35 [670]);
assign l_34[415]    = ( l_35 [671]);
assign l_34[416]    = ( l_35 [672]);
assign l_34[417]    = ( l_35 [673]);
assign l_34[418]    = ( l_35 [674]);
assign l_34[419]    = ( l_35 [675]);
assign l_34[420]    = ( l_35 [676]);
assign l_34[421]    = ( l_35 [677]);
assign l_34[422]    = ( l_35 [678]);
assign l_34[423]    = ( l_35 [679]);
assign l_34[424]    = ( l_35 [680]);
assign l_34[425]    = ( l_35 [681]);
assign l_34[426]    = ( l_35 [682]);
assign l_34[427]    = ( l_35 [683]);
assign l_34[428]    = ( l_35 [684]);
assign l_34[429]    = ( l_35 [685]);
assign l_34[430]    = ( l_35 [686]);
assign l_34[431]    = ( l_35 [687]);
assign l_34[432]    = ( l_35 [688]);
assign l_34[433]    = ( l_35 [689]);
assign l_34[434]    = ( l_35 [690]);
assign l_34[435]    = ( l_35 [691]);
assign l_34[436]    = ( l_35 [692]);
assign l_34[437]    = ( l_35 [693]);
assign l_34[438]    = ( l_35 [694]);
assign l_34[439]    = ( l_35 [695]);
assign l_34[440]    = ( l_35 [696]);
assign l_34[441]    = ( l_35 [697]);
assign l_34[442]    = ( l_35 [698]);
assign l_34[443]    = ( l_35 [699]);
assign l_34[444]    = ( l_35 [700]);
assign l_34[445]    = ( l_35 [701]);
assign l_34[446]    = ( l_35 [702]);
assign l_34[447]    = ( l_35 [703]);
assign l_34[448]    = ( l_35 [704]);
assign l_34[449]    = ( l_35 [705]);
assign l_34[450]    = ( l_35 [706]);
assign l_34[451]    = ( l_35 [707]);
assign l_34[452]    = ( l_35 [708]);
assign l_34[453]    = ( l_35 [709]);
assign l_34[454]    = ( l_35 [710]);
assign l_34[455]    = ( l_35 [711]);
assign l_34[456]    = ( l_35 [712]);
assign l_34[457]    = ( l_35 [713]);
assign l_34[458]    = ( l_35 [714]);
assign l_34[459]    = ( l_35 [715]);
assign l_34[460]    = ( l_35 [716]);
assign l_34[461]    = ( l_35 [717]);
assign l_34[462]    = ( l_35 [718]);
assign l_34[463]    = ( l_35 [719]);
assign l_34[464]    = ( l_35 [720]);
assign l_34[465]    = ( l_35 [721]);
assign l_34[466]    = ( l_35 [722]);
assign l_34[467]    = ( l_35 [723]);
assign l_34[468]    = ( l_35 [724]);
assign l_34[469]    = ( l_35 [725]);
assign l_34[470]    = ( l_35 [726]);
assign l_34[471]    = ( l_35 [727]);
assign l_34[472]    = ( l_35 [728]);
assign l_34[473]    = ( l_35 [729]);
assign l_34[474]    = ( l_35 [730]);
assign l_34[475]    = ( l_35 [731]);
assign l_34[476]    = ( l_35 [732]);
assign l_34[477]    = ( l_35 [733]);
assign l_34[478]    = ( l_35 [734]);
assign l_34[479]    = ( l_35 [735]);
assign l_34[480]    = ( l_35 [736]);
assign l_34[481]    = ( l_35 [737]);
assign l_34[482]    = ( l_35 [738]);
assign l_34[483]    = ( l_35 [739]);
assign l_34[484]    = ( l_35 [740]);
assign l_34[485]    = ( l_35 [741]);
assign l_34[486]    = ( l_35 [742]);
assign l_34[487]    = ( l_35 [743]);
assign l_34[488]    = ( l_35 [744]);
assign l_34[489]    = ( l_35 [745]);
assign l_34[490]    = ( l_35 [746]);
assign l_34[491]    = ( l_35 [747]);
assign l_34[492]    = ( l_35 [748]);
assign l_34[493]    = ( l_35 [749]);
assign l_34[494]    = ( l_35 [750]);
assign l_34[495]    = ( l_35 [751]);
assign l_34[496]    = ( l_35 [752]);
assign l_34[497]    = ( l_35 [753]);
assign l_34[498]    = ( l_35 [754]);
assign l_34[499]    = ( l_35 [755]);
assign l_34[500]    = ( l_35 [756]);
assign l_34[501]    = ( l_35 [757]);
assign l_34[502]    = ( l_35 [758]);
assign l_34[503]    = ( l_35 [759]);
assign l_34[504]    = ( l_35 [760]);
assign l_34[505]    = ( l_35 [761]);
assign l_34[506]    = ( l_35 [762]);
assign l_34[507]    = ( l_35 [763]);
assign l_34[508]    = ( l_35 [764]);
assign l_34[509]    = ( l_35 [765]);
assign l_34[510]    = ( l_35 [766]);
assign l_34[511]    = ( l_35 [767]);
assign l_34[512]    = ( l_35 [768]);
assign l_34[513]    = ( l_35 [769]);
assign l_34[514]    = ( l_35 [770]);
assign l_34[515]    = ( l_35 [771]);
assign l_34[516]    = ( l_35 [772]);
assign l_34[517]    = ( l_35 [773]);
assign l_34[518]    = ( l_35 [774]);
assign l_34[519]    = ( l_35 [775]);
assign l_34[520]    = ( l_35 [776]);
assign l_34[521]    = ( l_35 [777]);
assign l_34[522]    = ( l_35 [778]);
assign l_34[523]    = ( l_35 [779]);
assign l_34[524]    = ( l_35 [780]);
assign l_34[525]    = ( l_35 [781]);
assign l_34[526]    = ( l_35 [782]);
assign l_34[527]    = ( l_35 [783]);
assign l_34[528]    = ( l_35 [784]);
assign l_34[529]    = ( l_35 [785]);
assign l_35[0]    = ( l_36 [0]);
assign l_35[1]    = ( l_36 [1] & !i[1812]);
assign l_35[2]    = ( l_36 [2] & !i[1812]);
assign l_35[3]    = (!i[1812]) | ( l_36 [3] &  i[1812]);
assign l_35[4]    = (!i[1812]) | ( l_36 [4] &  i[1812]);
assign l_35[5]    = ( l_36 [5] & !i[1812]);
assign l_35[6]    = ( l_36 [6] & !i[1812]);
assign l_35[7]    = (!i[1812]) | ( l_36 [7] &  i[1812]);
assign l_35[8]    = (!i[1812]) | ( l_36 [8] &  i[1812]);
assign l_35[9]    = ( l_36 [9] & !i[1812]) | ( l_36 [10] &  i[1812]);
assign l_35[10]    = ( l_36 [10]);
assign l_35[11]    = ( l_36 [11] & !i[1812]) | ( l_36 [10] &  i[1812]);
assign l_35[12]    = ( l_36 [10] & !i[1812]) | ( l_36 [12] &  i[1812]);
assign l_35[13]    = ( l_36 [10] & !i[1812]) | ( l_36 [13] &  i[1812]);
assign l_35[14]    = ( l_36 [14] & !i[1812]) | ( l_36 [10] &  i[1812]);
assign l_35[15]    = ( l_36 [15] & !i[1812]) | ( l_36 [10] &  i[1812]);
assign l_35[16]    = ( l_36 [10] & !i[1812]) | ( l_36 [16] &  i[1812]);
assign l_35[17]    = ( l_36 [10] & !i[1812]) | ( l_36 [17] &  i[1812]);
assign l_35[18]    = ( l_36 [18]);
assign l_35[19]    = ( l_36 [19]);
assign l_35[20]    = ( l_36 [20]);
assign l_35[21]    = ( l_36 [21]);
assign l_35[22]    = ( l_36 [22]);
assign l_35[23]    = ( l_36 [23]);
assign l_35[24]    = ( l_36 [24]);
assign l_35[25]    = ( l_36 [25]);
assign l_35[26]    = ( l_36 [26]);
assign l_35[27]    = ( l_36 [27]);
assign l_35[28]    = ( l_36 [28]);
assign l_35[29]    = ( l_36 [29]);
assign l_35[30]    = ( l_36 [30]);
assign l_35[31]    = ( l_36 [31]);
assign l_35[32]    = ( l_36 [32]);
assign l_35[33]    = ( l_36 [33]);
assign l_35[34]    = ( l_36 [34]);
assign l_35[35]    = ( l_36 [35]);
assign l_35[36]    = ( l_36 [36]);
assign l_35[37]    = ( l_36 [37]);
assign l_35[38]    = ( l_36 [38]);
assign l_35[39]    = ( l_36 [39]);
assign l_35[40]    = ( l_36 [40]);
assign l_35[41]    = ( l_36 [41]);
assign l_35[42]    = ( l_36 [42]);
assign l_35[43]    = ( l_36 [43]);
assign l_35[44]    = ( l_36 [44]);
assign l_35[45]    = ( l_36 [45]);
assign l_35[46]    = ( l_36 [46]);
assign l_35[47]    = ( l_36 [47]);
assign l_35[48]    = ( l_36 [48]);
assign l_35[49]    = ( l_36 [49]);
assign l_35[50]    = ( l_36 [50]);
assign l_35[51]    = ( l_36 [51]);
assign l_35[52]    = ( l_36 [52]);
assign l_35[53]    = ( l_36 [53]);
assign l_35[54]    = ( l_36 [54]);
assign l_35[55]    = ( l_36 [55]);
assign l_35[56]    = ( l_36 [56]);
assign l_35[57]    = ( l_36 [57]);
assign l_35[58]    = ( l_36 [58]);
assign l_35[59]    = ( l_36 [59]);
assign l_35[60]    = ( l_36 [60]);
assign l_35[61]    = ( l_36 [61]);
assign l_35[62]    = ( l_36 [62]);
assign l_35[63]    = ( l_36 [63]);
assign l_35[64]    = ( l_36 [64]);
assign l_35[65]    = ( l_36 [65]);
assign l_35[66]    = ( l_36 [66]);
assign l_35[67]    = ( l_36 [67]);
assign l_35[68]    = ( l_36 [68]);
assign l_35[69]    = ( l_36 [69]);
assign l_35[70]    = ( l_36 [70]);
assign l_35[71]    = ( l_36 [71]);
assign l_35[72]    = ( l_36 [72]);
assign l_35[73]    = ( l_36 [73]);
assign l_35[74]    = ( l_36 [74]);
assign l_35[75]    = ( l_36 [75]);
assign l_35[76]    = ( l_36 [76]);
assign l_35[77]    = ( l_36 [77]);
assign l_35[78]    = ( l_36 [78]);
assign l_35[79]    = ( l_36 [79]);
assign l_35[80]    = ( l_36 [80]);
assign l_35[81]    = ( l_36 [81]);
assign l_35[82]    = ( l_36 [82]);
assign l_35[83]    = ( l_36 [83]);
assign l_35[84]    = ( l_36 [84]);
assign l_35[85]    = ( l_36 [85]);
assign l_35[86]    = ( l_36 [86]);
assign l_35[87]    = ( l_36 [87]);
assign l_35[88]    = ( l_36 [88]);
assign l_35[89]    = ( l_36 [89]);
assign l_35[90]    = ( l_36 [90]);
assign l_35[91]    = ( l_36 [91]);
assign l_35[92]    = ( l_36 [92]);
assign l_35[93]    = ( l_36 [93]);
assign l_35[94]    = ( l_36 [94]);
assign l_35[95]    = ( l_36 [95]);
assign l_35[96]    = ( l_36 [96]);
assign l_35[97]    = ( l_36 [97]);
assign l_35[98]    = ( l_36 [98]);
assign l_35[99]    = ( l_36 [99]);
assign l_35[100]    = ( l_36 [100]);
assign l_35[101]    = ( l_36 [101]);
assign l_35[102]    = ( l_36 [102]);
assign l_35[103]    = ( l_36 [103]);
assign l_35[104]    = ( l_36 [104]);
assign l_35[105]    = ( l_36 [105]);
assign l_35[106]    = ( l_36 [106]);
assign l_35[107]    = ( l_36 [107]);
assign l_35[108]    = ( l_36 [108]);
assign l_35[109]    = ( l_36 [109]);
assign l_35[110]    = ( l_36 [110]);
assign l_35[111]    = ( l_36 [111]);
assign l_35[112]    = ( l_36 [112]);
assign l_35[113]    = ( l_36 [113]);
assign l_35[114]    = ( l_36 [114]);
assign l_35[115]    = ( l_36 [115]);
assign l_35[116]    = ( l_36 [116]);
assign l_35[117]    = ( l_36 [117]);
assign l_35[118]    = ( l_36 [118]);
assign l_35[119]    = ( l_36 [119]);
assign l_35[120]    = ( l_36 [120]);
assign l_35[121]    = ( l_36 [121]);
assign l_35[122]    = ( l_36 [122]);
assign l_35[123]    = ( l_36 [123]);
assign l_35[124]    = ( l_36 [124]);
assign l_35[125]    = ( l_36 [125]);
assign l_35[126]    = ( l_36 [126]);
assign l_35[127]    = ( l_36 [127]);
assign l_35[128]    = ( l_36 [128]);
assign l_35[129]    = ( l_36 [129]);
assign l_35[130]    = ( l_36 [130]);
assign l_35[131]    = ( l_36 [131]);
assign l_35[132]    = ( l_36 [132]);
assign l_35[133]    = ( l_36 [133]);
assign l_35[134]    = ( l_36 [134]);
assign l_35[135]    = ( l_36 [135]);
assign l_35[136]    = ( l_36 [136]);
assign l_35[137]    = ( l_36 [137]);
assign l_35[138]    = ( l_36 [138]);
assign l_35[139]    = ( l_36 [139]);
assign l_35[140]    = ( l_36 [140]);
assign l_35[141]    = ( l_36 [141]);
assign l_35[142]    = ( l_36 [142]);
assign l_35[143]    = ( l_36 [143]);
assign l_35[144]    = ( l_36 [144]);
assign l_35[145]    = ( l_36 [145]);
assign l_35[146]    = ( l_36 [146]);
assign l_35[147]    = ( l_36 [147]);
assign l_35[148]    = ( l_36 [148]);
assign l_35[149]    = ( l_36 [149]);
assign l_35[150]    = ( l_36 [150]);
assign l_35[151]    = ( l_36 [151]);
assign l_35[152]    = ( l_36 [152]);
assign l_35[153]    = ( l_36 [153]);
assign l_35[154]    = ( l_36 [154]);
assign l_35[155]    = ( l_36 [155]);
assign l_35[156]    = ( l_36 [156]);
assign l_35[157]    = ( l_36 [157]);
assign l_35[158]    = ( l_36 [158]);
assign l_35[159]    = ( l_36 [159]);
assign l_35[160]    = ( l_36 [160]);
assign l_35[161]    = ( l_36 [161]);
assign l_35[162]    = ( l_36 [162]);
assign l_35[163]    = ( l_36 [163]);
assign l_35[164]    = ( l_36 [164]);
assign l_35[165]    = ( l_36 [165]);
assign l_35[166]    = ( l_36 [166]);
assign l_35[167]    = ( l_36 [167]);
assign l_35[168]    = ( l_36 [168]);
assign l_35[169]    = ( l_36 [169]);
assign l_35[170]    = ( l_36 [170]);
assign l_35[171]    = ( l_36 [171]);
assign l_35[172]    = ( l_36 [172]);
assign l_35[173]    = ( l_36 [173]);
assign l_35[174]    = ( l_36 [174]);
assign l_35[175]    = ( l_36 [175]);
assign l_35[176]    = ( l_36 [176]);
assign l_35[177]    = ( l_36 [177]);
assign l_35[178]    = ( l_36 [178]);
assign l_35[179]    = ( l_36 [179]);
assign l_35[180]    = ( l_36 [180]);
assign l_35[181]    = ( l_36 [181]);
assign l_35[182]    = ( l_36 [182]);
assign l_35[183]    = ( l_36 [183]);
assign l_35[184]    = ( l_36 [184]);
assign l_35[185]    = ( l_36 [185]);
assign l_35[186]    = ( l_36 [186]);
assign l_35[187]    = ( l_36 [187]);
assign l_35[188]    = ( l_36 [188]);
assign l_35[189]    = ( l_36 [189]);
assign l_35[190]    = ( l_36 [190]);
assign l_35[191]    = ( l_36 [191]);
assign l_35[192]    = ( l_36 [192]);
assign l_35[193]    = ( l_36 [193]);
assign l_35[194]    = ( l_36 [194]);
assign l_35[195]    = ( l_36 [195]);
assign l_35[196]    = ( l_36 [196]);
assign l_35[197]    = ( l_36 [197]);
assign l_35[198]    = ( l_36 [198]);
assign l_35[199]    = ( l_36 [199]);
assign l_35[200]    = ( l_36 [200]);
assign l_35[201]    = ( l_36 [201]);
assign l_35[202]    = ( l_36 [202]);
assign l_35[203]    = ( l_36 [203]);
assign l_35[204]    = ( l_36 [204]);
assign l_35[205]    = ( l_36 [205]);
assign l_35[206]    = ( l_36 [206]);
assign l_35[207]    = ( l_36 [207]);
assign l_35[208]    = ( l_36 [208]);
assign l_35[209]    = ( l_36 [209]);
assign l_35[210]    = ( l_36 [210]);
assign l_35[211]    = ( l_36 [211]);
assign l_35[212]    = ( l_36 [212]);
assign l_35[213]    = ( l_36 [213]);
assign l_35[214]    = ( l_36 [214]);
assign l_35[215]    = ( l_36 [215]);
assign l_35[216]    = ( l_36 [216]);
assign l_35[217]    = ( l_36 [217]);
assign l_35[218]    = ( l_36 [218]);
assign l_35[219]    = ( l_36 [219]);
assign l_35[220]    = ( l_36 [220]);
assign l_35[221]    = ( l_36 [221]);
assign l_35[222]    = ( l_36 [222]);
assign l_35[223]    = ( l_36 [223]);
assign l_35[224]    = ( l_36 [224]);
assign l_35[225]    = ( l_36 [225]);
assign l_35[226]    = ( l_36 [226]);
assign l_35[227]    = ( l_36 [227]);
assign l_35[228]    = ( l_36 [228]);
assign l_35[229]    = ( l_36 [229]);
assign l_35[230]    = ( l_36 [230]);
assign l_35[231]    = ( l_36 [231]);
assign l_35[232]    = ( l_36 [232]);
assign l_35[233]    = ( l_36 [233]);
assign l_35[234]    = ( l_36 [234]);
assign l_35[235]    = ( l_36 [235]);
assign l_35[236]    = ( l_36 [236]);
assign l_35[237]    = ( l_36 [237]);
assign l_35[238]    = ( l_36 [238]);
assign l_35[239]    = ( l_36 [239]);
assign l_35[240]    = ( l_36 [240]);
assign l_35[241]    = ( l_36 [241]);
assign l_35[242]    = ( l_36 [242]);
assign l_35[243]    = ( l_36 [243]);
assign l_35[244]    = ( l_36 [244]);
assign l_35[245]    = ( l_36 [245]);
assign l_35[246]    = ( l_36 [246]);
assign l_35[247]    = ( l_36 [247]);
assign l_35[248]    = ( l_36 [248]);
assign l_35[249]    = ( l_36 [249]);
assign l_35[250]    = ( l_36 [250]);
assign l_35[251]    = ( l_36 [251]);
assign l_35[252]    = ( l_36 [252]);
assign l_35[253]    = ( l_36 [253]);
assign l_35[254]    = ( l_36 [254]);
assign l_35[255]    = ( l_36 [255]);
assign l_35[256]    = ( l_36 [256]);
assign l_35[257]    = ( l_36 [257]);
assign l_35[258]    = ( l_36 [258]);
assign l_35[259]    = ( l_36 [259]);
assign l_35[260]    = ( l_36 [260]);
assign l_35[261]    = ( l_36 [261]);
assign l_35[262]    = ( l_36 [262]);
assign l_35[263]    = ( l_36 [263]);
assign l_35[264]    = ( l_36 [264]);
assign l_35[265]    = ( l_36 [265]);
assign l_35[266]    = ( l_36 [266]);
assign l_35[267]    = ( l_36 [267]);
assign l_35[268]    = ( l_36 [268]);
assign l_35[269]    = ( l_36 [269]);
assign l_35[270]    = ( l_36 [270]);
assign l_35[271]    = ( l_36 [271]);
assign l_35[272]    = ( l_36 [272]);
assign l_35[273]    = ( l_36 [273]);
assign l_35[274]    = ( l_36 [274]);
assign l_35[275]    = ( l_36 [275]);
assign l_35[276]    = ( l_36 [276]);
assign l_35[277]    = ( l_36 [277]);
assign l_35[278]    = ( l_36 [278]);
assign l_35[279]    = ( l_36 [279]);
assign l_35[280]    = ( l_36 [280]);
assign l_35[281]    = ( l_36 [281]);
assign l_35[282]    = ( l_36 [282]);
assign l_35[283]    = ( l_36 [283]);
assign l_35[284]    = ( l_36 [284]);
assign l_35[285]    = ( l_36 [285]);
assign l_35[286]    = ( l_36 [286]);
assign l_35[287]    = ( l_36 [287]);
assign l_35[288]    = ( l_36 [288]);
assign l_35[289]    = ( l_36 [289]);
assign l_35[290]    = ( l_36 [290]);
assign l_35[291]    = ( l_36 [291]);
assign l_35[292]    = ( l_36 [292]);
assign l_35[293]    = ( l_36 [293]);
assign l_35[294]    = ( l_36 [294]);
assign l_35[295]    = ( l_36 [295]);
assign l_35[296]    = ( l_36 [296]);
assign l_35[297]    = ( l_36 [297]);
assign l_35[298]    = ( l_36 [298]);
assign l_35[299]    = ( l_36 [299]);
assign l_35[300]    = ( l_36 [300]);
assign l_35[301]    = ( l_36 [301]);
assign l_35[302]    = ( l_36 [302]);
assign l_35[303]    = ( l_36 [303]);
assign l_35[304]    = ( l_36 [304]);
assign l_35[305]    = ( l_36 [305]);
assign l_35[306]    = ( l_36 [306]);
assign l_35[307]    = ( l_36 [307]);
assign l_35[308]    = ( l_36 [308]);
assign l_35[309]    = ( l_36 [309]);
assign l_35[310]    = ( l_36 [310]);
assign l_35[311]    = ( l_36 [311]);
assign l_35[312]    = ( l_36 [312]);
assign l_35[313]    = ( l_36 [313]);
assign l_35[314]    = ( l_36 [314]);
assign l_35[315]    = ( l_36 [315]);
assign l_35[316]    = ( l_36 [316]);
assign l_35[317]    = ( l_36 [317]);
assign l_35[318]    = ( l_36 [318]);
assign l_35[319]    = ( l_36 [319]);
assign l_35[320]    = ( l_36 [320]);
assign l_35[321]    = ( l_36 [321]);
assign l_35[322]    = ( l_36 [322]);
assign l_35[323]    = ( l_36 [323]);
assign l_35[324]    = ( l_36 [324]);
assign l_35[325]    = ( l_36 [325]);
assign l_35[326]    = ( l_36 [326]);
assign l_35[327]    = ( l_36 [327]);
assign l_35[328]    = ( l_36 [328]);
assign l_35[329]    = ( l_36 [329]);
assign l_35[330]    = ( l_36 [330]);
assign l_35[331]    = ( l_36 [331]);
assign l_35[332]    = ( l_36 [332]);
assign l_35[333]    = ( l_36 [333]);
assign l_35[334]    = ( l_36 [334]);
assign l_35[335]    = ( l_36 [335]);
assign l_35[336]    = ( l_36 [336]);
assign l_35[337]    = ( l_36 [337]);
assign l_35[338]    = ( l_36 [338]);
assign l_35[339]    = ( l_36 [339]);
assign l_35[340]    = ( l_36 [340]);
assign l_35[341]    = ( l_36 [341]);
assign l_35[342]    = ( l_36 [342]);
assign l_35[343]    = ( l_36 [343]);
assign l_35[344]    = ( l_36 [344]);
assign l_35[345]    = ( l_36 [345]);
assign l_35[346]    = ( l_36 [346]);
assign l_35[347]    = ( l_36 [347]);
assign l_35[348]    = ( l_36 [348]);
assign l_35[349]    = ( l_36 [349]);
assign l_35[350]    = ( l_36 [350]);
assign l_35[351]    = ( l_36 [351]);
assign l_35[352]    = ( l_36 [352]);
assign l_35[353]    = ( l_36 [353]);
assign l_35[354]    = ( l_36 [354]);
assign l_35[355]    = ( l_36 [355]);
assign l_35[356]    = ( l_36 [356]);
assign l_35[357]    = ( l_36 [357]);
assign l_35[358]    = ( l_36 [358]);
assign l_35[359]    = ( l_36 [359]);
assign l_35[360]    = ( l_36 [360]);
assign l_35[361]    = ( l_36 [361]);
assign l_35[362]    = ( l_36 [362]);
assign l_35[363]    = ( l_36 [363]);
assign l_35[364]    = ( l_36 [364]);
assign l_35[365]    = ( l_36 [365]);
assign l_35[366]    = ( l_36 [366]);
assign l_35[367]    = ( l_36 [367]);
assign l_35[368]    = ( l_36 [368]);
assign l_35[369]    = ( l_36 [369]);
assign l_35[370]    = ( l_36 [370]);
assign l_35[371]    = ( l_36 [371]);
assign l_35[372]    = ( l_36 [372]);
assign l_35[373]    = ( l_36 [373]);
assign l_35[374]    = ( l_36 [374]);
assign l_35[375]    = ( l_36 [375]);
assign l_35[376]    = ( l_36 [376]);
assign l_35[377]    = ( l_36 [377]);
assign l_35[378]    = ( l_36 [378]);
assign l_35[379]    = ( l_36 [379]);
assign l_35[380]    = ( l_36 [380]);
assign l_35[381]    = ( l_36 [381]);
assign l_35[382]    = ( l_36 [382]);
assign l_35[383]    = ( l_36 [383]);
assign l_35[384]    = ( l_36 [384]);
assign l_35[385]    = ( l_36 [385]);
assign l_35[386]    = ( l_36 [386]);
assign l_35[387]    = ( l_36 [387]);
assign l_35[388]    = ( l_36 [388]);
assign l_35[389]    = ( l_36 [389]);
assign l_35[390]    = ( l_36 [390]);
assign l_35[391]    = ( l_36 [391]);
assign l_35[392]    = ( l_36 [392]);
assign l_35[393]    = ( l_36 [393]);
assign l_35[394]    = ( l_36 [394]);
assign l_35[395]    = ( l_36 [395]);
assign l_35[396]    = ( l_36 [396]);
assign l_35[397]    = ( l_36 [397]);
assign l_35[398]    = ( l_36 [398]);
assign l_35[399]    = ( l_36 [399]);
assign l_35[400]    = ( l_36 [400]);
assign l_35[401]    = ( l_36 [401]);
assign l_35[402]    = ( l_36 [402]);
assign l_35[403]    = ( l_36 [403]);
assign l_35[404]    = ( l_36 [404]);
assign l_35[405]    = ( l_36 [405]);
assign l_35[406]    = ( l_36 [406]);
assign l_35[407]    = ( l_36 [407]);
assign l_35[408]    = ( l_36 [408]);
assign l_35[409]    = ( l_36 [409]);
assign l_35[410]    = ( l_36 [410]);
assign l_35[411]    = ( l_36 [411]);
assign l_35[412]    = ( l_36 [412]);
assign l_35[413]    = ( l_36 [413]);
assign l_35[414]    = ( l_36 [414]);
assign l_35[415]    = ( l_36 [415]);
assign l_35[416]    = ( l_36 [416]);
assign l_35[417]    = ( l_36 [417]);
assign l_35[418]    = ( l_36 [418]);
assign l_35[419]    = ( l_36 [419]);
assign l_35[420]    = ( l_36 [420]);
assign l_35[421]    = ( l_36 [421]);
assign l_35[422]    = ( l_36 [422]);
assign l_35[423]    = ( l_36 [423]);
assign l_35[424]    = ( l_36 [424]);
assign l_35[425]    = ( l_36 [425]);
assign l_35[426]    = ( l_36 [426]);
assign l_35[427]    = ( l_36 [427]);
assign l_35[428]    = ( l_36 [428]);
assign l_35[429]    = ( l_36 [429]);
assign l_35[430]    = ( l_36 [430]);
assign l_35[431]    = ( l_36 [431]);
assign l_35[432]    = ( l_36 [432]);
assign l_35[433]    = ( l_36 [433]);
assign l_35[434]    = ( l_36 [434]);
assign l_35[435]    = ( l_36 [435]);
assign l_35[436]    = ( l_36 [436]);
assign l_35[437]    = ( l_36 [437]);
assign l_35[438]    = ( l_36 [438]);
assign l_35[439]    = ( l_36 [439]);
assign l_35[440]    = ( l_36 [440]);
assign l_35[441]    = ( l_36 [441]);
assign l_35[442]    = ( l_36 [442]);
assign l_35[443]    = ( l_36 [443]);
assign l_35[444]    = ( l_36 [444]);
assign l_35[445]    = ( l_36 [445]);
assign l_35[446]    = ( l_36 [446]);
assign l_35[447]    = ( l_36 [447]);
assign l_35[448]    = ( l_36 [448]);
assign l_35[449]    = ( l_36 [449]);
assign l_35[450]    = ( l_36 [450]);
assign l_35[451]    = ( l_36 [451]);
assign l_35[452]    = ( l_36 [452]);
assign l_35[453]    = ( l_36 [453]);
assign l_35[454]    = ( l_36 [454]);
assign l_35[455]    = ( l_36 [455]);
assign l_35[456]    = ( l_36 [456]);
assign l_35[457]    = ( l_36 [457]);
assign l_35[458]    = ( l_36 [458]);
assign l_35[459]    = ( l_36 [459]);
assign l_35[460]    = ( l_36 [460]);
assign l_35[461]    = ( l_36 [461]);
assign l_35[462]    = ( l_36 [462]);
assign l_35[463]    = ( l_36 [463]);
assign l_35[464]    = ( l_36 [464]);
assign l_35[465]    = ( l_36 [465]);
assign l_35[466]    = ( l_36 [466]);
assign l_35[467]    = ( l_36 [467]);
assign l_35[468]    = ( l_36 [468]);
assign l_35[469]    = ( l_36 [469]);
assign l_35[470]    = ( l_36 [470]);
assign l_35[471]    = ( l_36 [471]);
assign l_35[472]    = ( l_36 [472]);
assign l_35[473]    = ( l_36 [473]);
assign l_35[474]    = ( l_36 [474]);
assign l_35[475]    = ( l_36 [475]);
assign l_35[476]    = ( l_36 [476]);
assign l_35[477]    = ( l_36 [477]);
assign l_35[478]    = ( l_36 [478]);
assign l_35[479]    = ( l_36 [479]);
assign l_35[480]    = ( l_36 [480]);
assign l_35[481]    = ( l_36 [481]);
assign l_35[482]    = ( l_36 [482]);
assign l_35[483]    = ( l_36 [483]);
assign l_35[484]    = ( l_36 [484]);
assign l_35[485]    = ( l_36 [485]);
assign l_35[486]    = ( l_36 [486]);
assign l_35[487]    = ( l_36 [487]);
assign l_35[488]    = ( l_36 [488]);
assign l_35[489]    = ( l_36 [489]);
assign l_35[490]    = ( l_36 [490]);
assign l_35[491]    = ( l_36 [491]);
assign l_35[492]    = ( l_36 [492]);
assign l_35[493]    = ( l_36 [493]);
assign l_35[494]    = ( l_36 [494]);
assign l_35[495]    = ( l_36 [495]);
assign l_35[496]    = ( l_36 [496]);
assign l_35[497]    = ( l_36 [497]);
assign l_35[498]    = ( l_36 [498]);
assign l_35[499]    = ( l_36 [499]);
assign l_35[500]    = ( l_36 [500]);
assign l_35[501]    = ( l_36 [501]);
assign l_35[502]    = ( l_36 [502]);
assign l_35[503]    = ( l_36 [503]);
assign l_35[504]    = ( l_36 [504]);
assign l_35[505]    = ( l_36 [505]);
assign l_35[506]    = ( l_36 [506]);
assign l_35[507]    = ( l_36 [507]);
assign l_35[508]    = ( l_36 [508]);
assign l_35[509]    = ( l_36 [509]);
assign l_35[510]    = ( l_36 [510]);
assign l_35[511]    = ( l_36 [511]);
assign l_35[512]    = ( l_36 [512]);
assign l_35[513]    = ( l_36 [513]);
assign l_35[514]    = ( l_36 [514]);
assign l_35[515]    = ( l_36 [515]);
assign l_35[516]    = ( l_36 [516]);
assign l_35[517]    = ( l_36 [517]);
assign l_35[518]    = ( l_36 [518]);
assign l_35[519]    = ( l_36 [519]);
assign l_35[520]    = ( l_36 [520]);
assign l_35[521]    = ( l_36 [521]);
assign l_35[522]    = ( l_36 [522]);
assign l_35[523]    = ( l_36 [523]);
assign l_35[524]    = ( l_36 [524]);
assign l_35[525]    = ( l_36 [525]);
assign l_35[526]    = ( l_36 [526]);
assign l_35[527]    = ( l_36 [527]);
assign l_35[528]    = ( l_36 [528]);
assign l_35[529]    = ( l_36 [529]);
assign l_35[530]    = ( l_36 [530] & !i[1812]) | ( l_36 [531] &  i[1812]);
assign l_35[531]    = ( l_36 [532] & !i[1812]) | ( l_36 [533] &  i[1812]);
assign l_35[532]    = ( l_36 [534] & !i[1812]) | ( l_36 [535] &  i[1812]);
assign l_35[533]    = ( l_36 [536] & !i[1812]) | ( l_36 [537] &  i[1812]);
assign l_35[534]    = ( l_36 [538] & !i[1812]) | ( l_36 [539] &  i[1812]);
assign l_35[535]    = ( l_36 [540] & !i[1812]) | ( l_36 [541] &  i[1812]);
assign l_35[536]    = ( l_36 [542] & !i[1812]) | ( l_36 [543] &  i[1812]);
assign l_35[537]    = ( l_36 [544] & !i[1812]) | ( l_36 [545] &  i[1812]);
assign l_35[538]    = ( l_36 [546] & !i[1812]) | ( l_36 [547] &  i[1812]);
assign l_35[539]    = ( l_36 [548] & !i[1812]) | ( l_36 [549] &  i[1812]);
assign l_35[540]    = ( l_36 [550] & !i[1812]) | ( l_36 [551] &  i[1812]);
assign l_35[541]    = ( l_36 [552] & !i[1812]) | ( l_36 [553] &  i[1812]);
assign l_35[542]    = ( l_36 [554] & !i[1812]) | ( l_36 [555] &  i[1812]);
assign l_35[543]    = ( l_36 [556] & !i[1812]) | ( l_36 [557] &  i[1812]);
assign l_35[544]    = ( l_36 [558] & !i[1812]) | ( l_36 [559] &  i[1812]);
assign l_35[545]    = ( l_36 [560] & !i[1812]) | ( l_36 [561] &  i[1812]);
assign l_35[546]    = ( l_36 [562] & !i[1812]) | ( l_36 [563] &  i[1812]);
assign l_35[547]    = ( l_36 [564] & !i[1812]) | ( l_36 [565] &  i[1812]);
assign l_35[548]    = ( l_36 [566] & !i[1812]) | ( l_36 [567] &  i[1812]);
assign l_35[549]    = ( l_36 [568] & !i[1812]) | ( l_36 [569] &  i[1812]);
assign l_35[550]    = ( l_36 [570] & !i[1812]) | ( l_36 [571] &  i[1812]);
assign l_35[551]    = ( l_36 [572] & !i[1812]) | ( l_36 [573] &  i[1812]);
assign l_35[552]    = ( l_36 [574] & !i[1812]) | ( l_36 [575] &  i[1812]);
assign l_35[553]    = ( l_36 [576] & !i[1812]) | ( l_36 [577] &  i[1812]);
assign l_35[554]    = ( l_36 [578] & !i[1812]) | ( l_36 [579] &  i[1812]);
assign l_35[555]    = ( l_36 [580] & !i[1812]) | ( l_36 [581] &  i[1812]);
assign l_35[556]    = ( l_36 [582] & !i[1812]) | ( l_36 [583] &  i[1812]);
assign l_35[557]    = ( l_36 [584] & !i[1812]) | ( l_36 [585] &  i[1812]);
assign l_35[558]    = ( l_36 [586] & !i[1812]) | ( l_36 [587] &  i[1812]);
assign l_35[559]    = ( l_36 [588] & !i[1812]) | ( l_36 [589] &  i[1812]);
assign l_35[560]    = ( l_36 [590] & !i[1812]) | ( l_36 [591] &  i[1812]);
assign l_35[561]    = ( l_36 [592] & !i[1812]) | ( l_36 [593] &  i[1812]);
assign l_35[562]    = ( l_36 [594] & !i[1812]) | ( l_36 [595] &  i[1812]);
assign l_35[563]    = ( l_36 [596] & !i[1812]) | ( l_36 [597] &  i[1812]);
assign l_35[564]    = ( l_36 [598] & !i[1812]) | ( l_36 [599] &  i[1812]);
assign l_35[565]    = ( l_36 [600] & !i[1812]) | ( l_36 [601] &  i[1812]);
assign l_35[566]    = ( l_36 [602] & !i[1812]) | ( l_36 [603] &  i[1812]);
assign l_35[567]    = ( l_36 [604] & !i[1812]) | ( l_36 [605] &  i[1812]);
assign l_35[568]    = ( l_36 [606] & !i[1812]) | ( l_36 [607] &  i[1812]);
assign l_35[569]    = ( l_36 [608] & !i[1812]) | ( l_36 [609] &  i[1812]);
assign l_35[570]    = ( l_36 [610] & !i[1812]) | ( l_36 [611] &  i[1812]);
assign l_35[571]    = ( l_36 [612] & !i[1812]) | ( l_36 [613] &  i[1812]);
assign l_35[572]    = ( l_36 [614] & !i[1812]) | ( l_36 [615] &  i[1812]);
assign l_35[573]    = ( l_36 [616] & !i[1812]) | ( l_36 [617] &  i[1812]);
assign l_35[574]    = ( l_36 [618] & !i[1812]) | ( l_36 [619] &  i[1812]);
assign l_35[575]    = ( l_36 [620] & !i[1812]) | ( l_36 [621] &  i[1812]);
assign l_35[576]    = ( l_36 [622] & !i[1812]) | ( l_36 [623] &  i[1812]);
assign l_35[577]    = ( l_36 [624] & !i[1812]) | ( l_36 [625] &  i[1812]);
assign l_35[578]    = ( l_36 [626] & !i[1812]) | ( l_36 [627] &  i[1812]);
assign l_35[579]    = ( l_36 [628] & !i[1812]) | ( l_36 [629] &  i[1812]);
assign l_35[580]    = ( l_36 [630] & !i[1812]) | ( l_36 [631] &  i[1812]);
assign l_35[581]    = ( l_36 [632] & !i[1812]) | ( l_36 [633] &  i[1812]);
assign l_35[582]    = ( l_36 [634] & !i[1812]) | ( l_36 [635] &  i[1812]);
assign l_35[583]    = ( l_36 [636] & !i[1812]) | ( l_36 [637] &  i[1812]);
assign l_35[584]    = ( l_36 [638] & !i[1812]) | ( l_36 [639] &  i[1812]);
assign l_35[585]    = ( l_36 [640] & !i[1812]) | ( l_36 [641] &  i[1812]);
assign l_35[586]    = ( l_36 [642] & !i[1812]) | ( l_36 [643] &  i[1812]);
assign l_35[587]    = ( l_36 [644] & !i[1812]) | ( l_36 [645] &  i[1812]);
assign l_35[588]    = ( l_36 [646] & !i[1812]) | ( l_36 [647] &  i[1812]);
assign l_35[589]    = ( l_36 [648] & !i[1812]) | ( l_36 [649] &  i[1812]);
assign l_35[590]    = ( l_36 [650] & !i[1812]) | ( l_36 [651] &  i[1812]);
assign l_35[591]    = ( l_36 [652] & !i[1812]) | ( l_36 [653] &  i[1812]);
assign l_35[592]    = ( l_36 [654] & !i[1812]) | ( l_36 [655] &  i[1812]);
assign l_35[593]    = ( l_36 [656] & !i[1812]) | ( l_36 [657] &  i[1812]);
assign l_35[594]    = ( l_36 [658] & !i[1812]) | ( l_36 [659] &  i[1812]);
assign l_35[595]    = ( l_36 [660] & !i[1812]) | ( l_36 [661] &  i[1812]);
assign l_35[596]    = ( l_36 [662] & !i[1812]) | ( l_36 [663] &  i[1812]);
assign l_35[597]    = ( l_36 [664] & !i[1812]) | ( l_36 [665] &  i[1812]);
assign l_35[598]    = ( l_36 [666] & !i[1812]) | ( l_36 [667] &  i[1812]);
assign l_35[599]    = ( l_36 [668] & !i[1812]) | ( l_36 [669] &  i[1812]);
assign l_35[600]    = ( l_36 [670] & !i[1812]) | ( l_36 [671] &  i[1812]);
assign l_35[601]    = ( l_36 [672] & !i[1812]) | ( l_36 [673] &  i[1812]);
assign l_35[602]    = ( l_36 [674] & !i[1812]) | ( l_36 [675] &  i[1812]);
assign l_35[603]    = ( l_36 [676] & !i[1812]) | ( l_36 [677] &  i[1812]);
assign l_35[604]    = ( l_36 [678] & !i[1812]) | ( l_36 [679] &  i[1812]);
assign l_35[605]    = ( l_36 [680] & !i[1812]) | ( l_36 [681] &  i[1812]);
assign l_35[606]    = ( l_36 [682] & !i[1812]) | ( l_36 [683] &  i[1812]);
assign l_35[607]    = ( l_36 [684] & !i[1812]) | ( l_36 [685] &  i[1812]);
assign l_35[608]    = ( l_36 [686] & !i[1812]) | ( l_36 [687] &  i[1812]);
assign l_35[609]    = ( l_36 [688] & !i[1812]) | ( l_36 [689] &  i[1812]);
assign l_35[610]    = ( l_36 [690] & !i[1812]) | ( l_36 [691] &  i[1812]);
assign l_35[611]    = ( l_36 [692] & !i[1812]) | ( l_36 [693] &  i[1812]);
assign l_35[612]    = ( l_36 [694] & !i[1812]) | ( l_36 [695] &  i[1812]);
assign l_35[613]    = ( l_36 [696] & !i[1812]) | ( l_36 [697] &  i[1812]);
assign l_35[614]    = ( l_36 [698] & !i[1812]) | ( l_36 [699] &  i[1812]);
assign l_35[615]    = ( l_36 [700] & !i[1812]) | ( l_36 [701] &  i[1812]);
assign l_35[616]    = ( l_36 [702] & !i[1812]) | ( l_36 [703] &  i[1812]);
assign l_35[617]    = ( l_36 [704] & !i[1812]) | ( l_36 [705] &  i[1812]);
assign l_35[618]    = ( l_36 [706] & !i[1812]) | ( l_36 [707] &  i[1812]);
assign l_35[619]    = ( l_36 [708] & !i[1812]) | ( l_36 [709] &  i[1812]);
assign l_35[620]    = ( l_36 [710] & !i[1812]) | ( l_36 [711] &  i[1812]);
assign l_35[621]    = ( l_36 [712] & !i[1812]) | ( l_36 [713] &  i[1812]);
assign l_35[622]    = ( l_36 [714] & !i[1812]) | ( l_36 [715] &  i[1812]);
assign l_35[623]    = ( l_36 [716] & !i[1812]) | ( l_36 [717] &  i[1812]);
assign l_35[624]    = ( l_36 [718] & !i[1812]) | ( l_36 [719] &  i[1812]);
assign l_35[625]    = ( l_36 [720] & !i[1812]) | ( l_36 [721] &  i[1812]);
assign l_35[626]    = ( l_36 [722] & !i[1812]) | ( l_36 [723] &  i[1812]);
assign l_35[627]    = ( l_36 [724] & !i[1812]) | ( l_36 [725] &  i[1812]);
assign l_35[628]    = ( l_36 [726] & !i[1812]) | ( l_36 [727] &  i[1812]);
assign l_35[629]    = ( l_36 [728] & !i[1812]) | ( l_36 [729] &  i[1812]);
assign l_35[630]    = ( l_36 [730] & !i[1812]) | ( l_36 [731] &  i[1812]);
assign l_35[631]    = ( l_36 [732] & !i[1812]) | ( l_36 [733] &  i[1812]);
assign l_35[632]    = ( l_36 [734] & !i[1812]) | ( l_36 [735] &  i[1812]);
assign l_35[633]    = ( l_36 [736] & !i[1812]) | ( l_36 [737] &  i[1812]);
assign l_35[634]    = ( l_36 [738] & !i[1812]) | ( l_36 [739] &  i[1812]);
assign l_35[635]    = ( l_36 [740] & !i[1812]) | ( l_36 [741] &  i[1812]);
assign l_35[636]    = ( l_36 [742] & !i[1812]) | ( l_36 [743] &  i[1812]);
assign l_35[637]    = ( l_36 [744] & !i[1812]) | ( l_36 [745] &  i[1812]);
assign l_35[638]    = ( l_36 [746] & !i[1812]) | ( l_36 [747] &  i[1812]);
assign l_35[639]    = ( l_36 [748] & !i[1812]) | ( l_36 [749] &  i[1812]);
assign l_35[640]    = ( l_36 [750] & !i[1812]) | ( l_36 [751] &  i[1812]);
assign l_35[641]    = ( l_36 [752] & !i[1812]) | ( l_36 [753] &  i[1812]);
assign l_35[642]    = ( l_36 [754] & !i[1812]) | ( l_36 [755] &  i[1812]);
assign l_35[643]    = ( l_36 [756] & !i[1812]) | ( l_36 [757] &  i[1812]);
assign l_35[644]    = ( l_36 [758] & !i[1812]) | ( l_36 [759] &  i[1812]);
assign l_35[645]    = ( l_36 [760] & !i[1812]) | ( l_36 [761] &  i[1812]);
assign l_35[646]    = ( l_36 [762] & !i[1812]) | ( l_36 [763] &  i[1812]);
assign l_35[647]    = ( l_36 [764] & !i[1812]) | ( l_36 [765] &  i[1812]);
assign l_35[648]    = ( l_36 [766] & !i[1812]) | ( l_36 [767] &  i[1812]);
assign l_35[649]    = ( l_36 [768] & !i[1812]) | ( l_36 [769] &  i[1812]);
assign l_35[650]    = ( l_36 [770] & !i[1812]) | ( l_36 [771] &  i[1812]);
assign l_35[651]    = ( l_36 [772] & !i[1812]) | ( l_36 [773] &  i[1812]);
assign l_35[652]    = ( l_36 [774] & !i[1812]) | ( l_36 [775] &  i[1812]);
assign l_35[653]    = ( l_36 [776] & !i[1812]) | ( l_36 [777] &  i[1812]);
assign l_35[654]    = ( l_36 [778] & !i[1812]) | ( l_36 [779] &  i[1812]);
assign l_35[655]    = ( l_36 [780] & !i[1812]) | ( l_36 [781] &  i[1812]);
assign l_35[656]    = ( l_36 [782] & !i[1812]) | ( l_36 [783] &  i[1812]);
assign l_35[657]    = ( l_36 [784] & !i[1812]) | ( l_36 [785] &  i[1812]);
assign l_35[658]    = ( l_36 [786] & !i[1812]) | ( l_36 [787] &  i[1812]);
assign l_35[659]    = ( l_36 [788] & !i[1812]) | ( l_36 [789] &  i[1812]);
assign l_35[660]    = ( l_36 [790] & !i[1812]) | ( l_36 [791] &  i[1812]);
assign l_35[661]    = ( l_36 [792] & !i[1812]) | ( l_36 [793] &  i[1812]);
assign l_35[662]    = ( l_36 [794] & !i[1812]) | ( l_36 [795] &  i[1812]);
assign l_35[663]    = ( l_36 [796] & !i[1812]) | ( l_36 [797] &  i[1812]);
assign l_35[664]    = ( l_36 [798] & !i[1812]) | ( l_36 [799] &  i[1812]);
assign l_35[665]    = ( l_36 [800] & !i[1812]) | ( l_36 [801] &  i[1812]);
assign l_35[666]    = ( l_36 [802] & !i[1812]) | ( l_36 [803] &  i[1812]);
assign l_35[667]    = ( l_36 [804] & !i[1812]) | ( l_36 [805] &  i[1812]);
assign l_35[668]    = ( l_36 [806] & !i[1812]) | ( l_36 [807] &  i[1812]);
assign l_35[669]    = ( l_36 [808] & !i[1812]) | ( l_36 [809] &  i[1812]);
assign l_35[670]    = ( l_36 [810] & !i[1812]) | ( l_36 [811] &  i[1812]);
assign l_35[671]    = ( l_36 [812] & !i[1812]) | ( l_36 [813] &  i[1812]);
assign l_35[672]    = ( l_36 [814] & !i[1812]) | ( l_36 [815] &  i[1812]);
assign l_35[673]    = ( l_36 [816] & !i[1812]) | ( l_36 [817] &  i[1812]);
assign l_35[674]    = ( l_36 [818] & !i[1812]) | ( l_36 [819] &  i[1812]);
assign l_35[675]    = ( l_36 [820] & !i[1812]) | ( l_36 [821] &  i[1812]);
assign l_35[676]    = ( l_36 [822] & !i[1812]) | ( l_36 [823] &  i[1812]);
assign l_35[677]    = ( l_36 [824] & !i[1812]) | ( l_36 [825] &  i[1812]);
assign l_35[678]    = ( l_36 [826] & !i[1812]) | ( l_36 [827] &  i[1812]);
assign l_35[679]    = ( l_36 [828] & !i[1812]) | ( l_36 [829] &  i[1812]);
assign l_35[680]    = ( l_36 [830] & !i[1812]) | ( l_36 [831] &  i[1812]);
assign l_35[681]    = ( l_36 [832] & !i[1812]) | ( l_36 [833] &  i[1812]);
assign l_35[682]    = ( l_36 [834] & !i[1812]) | ( l_36 [835] &  i[1812]);
assign l_35[683]    = ( l_36 [836] & !i[1812]) | ( l_36 [837] &  i[1812]);
assign l_35[684]    = ( l_36 [838] & !i[1812]) | ( l_36 [839] &  i[1812]);
assign l_35[685]    = ( l_36 [840] & !i[1812]) | ( l_36 [841] &  i[1812]);
assign l_35[686]    = ( l_36 [842] & !i[1812]) | ( l_36 [843] &  i[1812]);
assign l_35[687]    = ( l_36 [844] & !i[1812]) | ( l_36 [845] &  i[1812]);
assign l_35[688]    = ( l_36 [846] & !i[1812]) | ( l_36 [847] &  i[1812]);
assign l_35[689]    = ( l_36 [848] & !i[1812]) | ( l_36 [849] &  i[1812]);
assign l_35[690]    = ( l_36 [850] & !i[1812]) | ( l_36 [851] &  i[1812]);
assign l_35[691]    = ( l_36 [852] & !i[1812]) | ( l_36 [853] &  i[1812]);
assign l_35[692]    = ( l_36 [854] & !i[1812]) | ( l_36 [855] &  i[1812]);
assign l_35[693]    = ( l_36 [856] & !i[1812]) | ( l_36 [857] &  i[1812]);
assign l_35[694]    = ( l_36 [858] & !i[1812]) | ( l_36 [859] &  i[1812]);
assign l_35[695]    = ( l_36 [860] & !i[1812]) | ( l_36 [861] &  i[1812]);
assign l_35[696]    = ( l_36 [862] & !i[1812]) | ( l_36 [863] &  i[1812]);
assign l_35[697]    = ( l_36 [864] & !i[1812]) | ( l_36 [865] &  i[1812]);
assign l_35[698]    = ( l_36 [866] & !i[1812]) | ( l_36 [867] &  i[1812]);
assign l_35[699]    = ( l_36 [868] & !i[1812]) | ( l_36 [869] &  i[1812]);
assign l_35[700]    = ( l_36 [870] & !i[1812]) | ( l_36 [871] &  i[1812]);
assign l_35[701]    = ( l_36 [872] & !i[1812]) | ( l_36 [873] &  i[1812]);
assign l_35[702]    = ( l_36 [874] & !i[1812]) | ( l_36 [875] &  i[1812]);
assign l_35[703]    = ( l_36 [876] & !i[1812]) | ( l_36 [877] &  i[1812]);
assign l_35[704]    = ( l_36 [878] & !i[1812]) | ( l_36 [879] &  i[1812]);
assign l_35[705]    = ( l_36 [880] & !i[1812]) | ( l_36 [881] &  i[1812]);
assign l_35[706]    = ( l_36 [882] & !i[1812]) | ( l_36 [883] &  i[1812]);
assign l_35[707]    = ( l_36 [884] & !i[1812]) | ( l_36 [885] &  i[1812]);
assign l_35[708]    = ( l_36 [886] & !i[1812]) | ( l_36 [887] &  i[1812]);
assign l_35[709]    = ( l_36 [888] & !i[1812]) | ( l_36 [889] &  i[1812]);
assign l_35[710]    = ( l_36 [890] & !i[1812]) | ( l_36 [891] &  i[1812]);
assign l_35[711]    = ( l_36 [892] & !i[1812]) | ( l_36 [893] &  i[1812]);
assign l_35[712]    = ( l_36 [894] & !i[1812]) | ( l_36 [895] &  i[1812]);
assign l_35[713]    = ( l_36 [896] & !i[1812]) | ( l_36 [897] &  i[1812]);
assign l_35[714]    = ( l_36 [898] & !i[1812]) | ( l_36 [899] &  i[1812]);
assign l_35[715]    = ( l_36 [900] & !i[1812]) | ( l_36 [901] &  i[1812]);
assign l_35[716]    = ( l_36 [902] & !i[1812]) | ( l_36 [903] &  i[1812]);
assign l_35[717]    = ( l_36 [904] & !i[1812]) | ( l_36 [905] &  i[1812]);
assign l_35[718]    = ( l_36 [906] & !i[1812]) | ( l_36 [907] &  i[1812]);
assign l_35[719]    = ( l_36 [908] & !i[1812]) | ( l_36 [909] &  i[1812]);
assign l_35[720]    = ( l_36 [910] & !i[1812]) | ( l_36 [911] &  i[1812]);
assign l_35[721]    = ( l_36 [912] & !i[1812]) | ( l_36 [913] &  i[1812]);
assign l_35[722]    = ( l_36 [914] & !i[1812]) | ( l_36 [915] &  i[1812]);
assign l_35[723]    = ( l_36 [916] & !i[1812]) | ( l_36 [917] &  i[1812]);
assign l_35[724]    = ( l_36 [918] & !i[1812]) | ( l_36 [919] &  i[1812]);
assign l_35[725]    = ( l_36 [920] & !i[1812]) | ( l_36 [921] &  i[1812]);
assign l_35[726]    = ( l_36 [922] & !i[1812]) | ( l_36 [923] &  i[1812]);
assign l_35[727]    = ( l_36 [924] & !i[1812]) | ( l_36 [925] &  i[1812]);
assign l_35[728]    = ( l_36 [926] & !i[1812]) | ( l_36 [927] &  i[1812]);
assign l_35[729]    = ( l_36 [928] & !i[1812]) | ( l_36 [929] &  i[1812]);
assign l_35[730]    = ( l_36 [930] & !i[1812]) | ( l_36 [931] &  i[1812]);
assign l_35[731]    = ( l_36 [932] & !i[1812]) | ( l_36 [933] &  i[1812]);
assign l_35[732]    = ( l_36 [934] & !i[1812]) | ( l_36 [935] &  i[1812]);
assign l_35[733]    = ( l_36 [936] & !i[1812]) | ( l_36 [937] &  i[1812]);
assign l_35[734]    = ( l_36 [938] & !i[1812]) | ( l_36 [939] &  i[1812]);
assign l_35[735]    = ( l_36 [940] & !i[1812]) | ( l_36 [941] &  i[1812]);
assign l_35[736]    = ( l_36 [942] & !i[1812]) | ( l_36 [943] &  i[1812]);
assign l_35[737]    = ( l_36 [944] & !i[1812]) | ( l_36 [945] &  i[1812]);
assign l_35[738]    = ( l_36 [946] & !i[1812]) | ( l_36 [947] &  i[1812]);
assign l_35[739]    = ( l_36 [948] & !i[1812]) | ( l_36 [949] &  i[1812]);
assign l_35[740]    = ( l_36 [950] & !i[1812]) | ( l_36 [951] &  i[1812]);
assign l_35[741]    = ( l_36 [952] & !i[1812]) | ( l_36 [953] &  i[1812]);
assign l_35[742]    = ( l_36 [954] & !i[1812]) | ( l_36 [955] &  i[1812]);
assign l_35[743]    = ( l_36 [956] & !i[1812]) | ( l_36 [957] &  i[1812]);
assign l_35[744]    = ( l_36 [958] & !i[1812]) | ( l_36 [959] &  i[1812]);
assign l_35[745]    = ( l_36 [960] & !i[1812]) | ( l_36 [961] &  i[1812]);
assign l_35[746]    = ( l_36 [962] & !i[1812]) | ( l_36 [963] &  i[1812]);
assign l_35[747]    = ( l_36 [964] & !i[1812]) | ( l_36 [965] &  i[1812]);
assign l_35[748]    = ( l_36 [966] & !i[1812]) | ( l_36 [967] &  i[1812]);
assign l_35[749]    = ( l_36 [968] & !i[1812]) | ( l_36 [969] &  i[1812]);
assign l_35[750]    = ( l_36 [970] & !i[1812]) | ( l_36 [971] &  i[1812]);
assign l_35[751]    = ( l_36 [972] & !i[1812]) | ( l_36 [973] &  i[1812]);
assign l_35[752]    = ( l_36 [974] & !i[1812]) | ( l_36 [975] &  i[1812]);
assign l_35[753]    = ( l_36 [976] & !i[1812]) | ( l_36 [977] &  i[1812]);
assign l_35[754]    = ( l_36 [978] & !i[1812]) | ( l_36 [979] &  i[1812]);
assign l_35[755]    = ( l_36 [980] & !i[1812]) | ( l_36 [981] &  i[1812]);
assign l_35[756]    = ( l_36 [982] & !i[1812]) | ( l_36 [983] &  i[1812]);
assign l_35[757]    = ( l_36 [984] & !i[1812]) | ( l_36 [985] &  i[1812]);
assign l_35[758]    = ( l_36 [986] & !i[1812]) | ( l_36 [987] &  i[1812]);
assign l_35[759]    = ( l_36 [988] & !i[1812]) | ( l_36 [989] &  i[1812]);
assign l_35[760]    = ( l_36 [990] & !i[1812]) | ( l_36 [991] &  i[1812]);
assign l_35[761]    = ( l_36 [992] & !i[1812]) | ( l_36 [993] &  i[1812]);
assign l_35[762]    = ( l_36 [994] & !i[1812]) | ( l_36 [995] &  i[1812]);
assign l_35[763]    = ( l_36 [996] & !i[1812]) | ( l_36 [997] &  i[1812]);
assign l_35[764]    = ( l_36 [998] & !i[1812]) | ( l_36 [999] &  i[1812]);
assign l_35[765]    = ( l_36 [1000] & !i[1812]) | ( l_36 [1001] &  i[1812]);
assign l_35[766]    = ( l_36 [1002] & !i[1812]) | ( l_36 [1003] &  i[1812]);
assign l_35[767]    = ( l_36 [1004] & !i[1812]) | ( l_36 [1005] &  i[1812]);
assign l_35[768]    = ( l_36 [1006] & !i[1812]) | ( l_36 [1007] &  i[1812]);
assign l_35[769]    = ( l_36 [1008] & !i[1812]) | ( l_36 [1009] &  i[1812]);
assign l_35[770]    = ( l_36 [1010] & !i[1812]) | ( l_36 [1011] &  i[1812]);
assign l_35[771]    = ( l_36 [1012] & !i[1812]) | ( l_36 [1013] &  i[1812]);
assign l_35[772]    = ( l_36 [1014] & !i[1812]) | ( l_36 [1015] &  i[1812]);
assign l_35[773]    = ( l_36 [1016] & !i[1812]) | ( l_36 [1017] &  i[1812]);
assign l_35[774]    = ( l_36 [1018] & !i[1812]) | ( l_36 [1019] &  i[1812]);
assign l_35[775]    = ( l_36 [1020] & !i[1812]) | ( l_36 [1021] &  i[1812]);
assign l_35[776]    = ( l_36 [1022] & !i[1812]) | ( l_36 [1023] &  i[1812]);
assign l_35[777]    = ( l_36 [1024] & !i[1812]) | ( l_36 [1025] &  i[1812]);
assign l_35[778]    = ( l_36 [1026] & !i[1812]) | ( l_36 [1027] &  i[1812]);
assign l_35[779]    = ( l_36 [1028] & !i[1812]) | ( l_36 [1029] &  i[1812]);
assign l_35[780]    = ( l_36 [1030] & !i[1812]) | ( l_36 [1031] &  i[1812]);
assign l_35[781]    = ( l_36 [1032] & !i[1812]) | ( l_36 [1033] &  i[1812]);
assign l_35[782]    = ( l_36 [1034] & !i[1812]) | ( l_36 [1035] &  i[1812]);
assign l_35[783]    = ( l_36 [1036] & !i[1812]) | ( l_36 [1037] &  i[1812]);
assign l_35[784]    = ( l_36 [1038] & !i[1812]) | ( l_36 [1039] &  i[1812]);
assign l_35[785]    = ( l_36 [1040] & !i[1812]) | ( l_36 [1041] &  i[1812]);
assign l_36[0]    = ( l_37 [0]);
assign l_36[1]    = ( l_37 [1] & !i[1800]);
assign l_36[2]    = ( l_37 [2] & !i[1800]);
assign l_36[3]    = (!i[1800]) | ( l_37 [3] &  i[1800]);
assign l_36[4]    = (!i[1800]) | ( l_37 [4] &  i[1800]);
assign l_36[5]    = ( l_37 [5] & !i[1800]);
assign l_36[6]    = ( l_37 [6] & !i[1800]);
assign l_36[7]    = (!i[1800]) | ( l_37 [7] &  i[1800]);
assign l_36[8]    = (!i[1800]) | ( l_37 [8] &  i[1800]);
assign l_36[9]    = ( l_37 [9] & !i[1800]) | ( l_37 [10] &  i[1800]);
assign l_36[10]    = ( l_37 [10]);
assign l_36[11]    = ( l_37 [11] & !i[1800]) | ( l_37 [10] &  i[1800]);
assign l_36[12]    = ( l_37 [10] & !i[1800]) | ( l_37 [12] &  i[1800]);
assign l_36[13]    = ( l_37 [10] & !i[1800]) | ( l_37 [13] &  i[1800]);
assign l_36[14]    = ( l_37 [14] & !i[1800]) | ( l_37 [10] &  i[1800]);
assign l_36[15]    = ( l_37 [15] & !i[1800]) | ( l_37 [10] &  i[1800]);
assign l_36[16]    = ( l_37 [10] & !i[1800]) | ( l_37 [16] &  i[1800]);
assign l_36[17]    = ( l_37 [10] & !i[1800]) | ( l_37 [17] &  i[1800]);
assign l_36[18]    = ( l_37 [18]);
assign l_36[19]    = ( l_37 [19]);
assign l_36[20]    = ( l_37 [20]);
assign l_36[21]    = ( l_37 [21]);
assign l_36[22]    = ( l_37 [22]);
assign l_36[23]    = ( l_37 [23]);
assign l_36[24]    = ( l_37 [24]);
assign l_36[25]    = ( l_37 [25]);
assign l_36[26]    = ( l_37 [26]);
assign l_36[27]    = ( l_37 [27]);
assign l_36[28]    = ( l_37 [28]);
assign l_36[29]    = ( l_37 [29]);
assign l_36[30]    = ( l_37 [30]);
assign l_36[31]    = ( l_37 [31]);
assign l_36[32]    = ( l_37 [32]);
assign l_36[33]    = ( l_37 [33]);
assign l_36[34]    = ( l_37 [34]);
assign l_36[35]    = ( l_37 [35]);
assign l_36[36]    = ( l_37 [36]);
assign l_36[37]    = ( l_37 [37]);
assign l_36[38]    = ( l_37 [38]);
assign l_36[39]    = ( l_37 [39]);
assign l_36[40]    = ( l_37 [40]);
assign l_36[41]    = ( l_37 [41]);
assign l_36[42]    = ( l_37 [42]);
assign l_36[43]    = ( l_37 [43]);
assign l_36[44]    = ( l_37 [44]);
assign l_36[45]    = ( l_37 [45]);
assign l_36[46]    = ( l_37 [46]);
assign l_36[47]    = ( l_37 [47]);
assign l_36[48]    = ( l_37 [48]);
assign l_36[49]    = ( l_37 [49]);
assign l_36[50]    = ( l_37 [50]);
assign l_36[51]    = ( l_37 [51]);
assign l_36[52]    = ( l_37 [52]);
assign l_36[53]    = ( l_37 [53]);
assign l_36[54]    = ( l_37 [54]);
assign l_36[55]    = ( l_37 [55]);
assign l_36[56]    = ( l_37 [56]);
assign l_36[57]    = ( l_37 [57]);
assign l_36[58]    = ( l_37 [58]);
assign l_36[59]    = ( l_37 [59]);
assign l_36[60]    = ( l_37 [60]);
assign l_36[61]    = ( l_37 [61]);
assign l_36[62]    = ( l_37 [62]);
assign l_36[63]    = ( l_37 [63]);
assign l_36[64]    = ( l_37 [64]);
assign l_36[65]    = ( l_37 [65]);
assign l_36[66]    = ( l_37 [66]);
assign l_36[67]    = ( l_37 [67]);
assign l_36[68]    = ( l_37 [68]);
assign l_36[69]    = ( l_37 [69]);
assign l_36[70]    = ( l_37 [70]);
assign l_36[71]    = ( l_37 [71]);
assign l_36[72]    = ( l_37 [72]);
assign l_36[73]    = ( l_37 [73]);
assign l_36[74]    = ( l_37 [74]);
assign l_36[75]    = ( l_37 [75]);
assign l_36[76]    = ( l_37 [76]);
assign l_36[77]    = ( l_37 [77]);
assign l_36[78]    = ( l_37 [78]);
assign l_36[79]    = ( l_37 [79]);
assign l_36[80]    = ( l_37 [80]);
assign l_36[81]    = ( l_37 [81]);
assign l_36[82]    = ( l_37 [82]);
assign l_36[83]    = ( l_37 [83]);
assign l_36[84]    = ( l_37 [84]);
assign l_36[85]    = ( l_37 [85]);
assign l_36[86]    = ( l_37 [86]);
assign l_36[87]    = ( l_37 [87]);
assign l_36[88]    = ( l_37 [88]);
assign l_36[89]    = ( l_37 [89]);
assign l_36[90]    = ( l_37 [90]);
assign l_36[91]    = ( l_37 [91]);
assign l_36[92]    = ( l_37 [92]);
assign l_36[93]    = ( l_37 [93]);
assign l_36[94]    = ( l_37 [94]);
assign l_36[95]    = ( l_37 [95]);
assign l_36[96]    = ( l_37 [96]);
assign l_36[97]    = ( l_37 [97]);
assign l_36[98]    = ( l_37 [98]);
assign l_36[99]    = ( l_37 [99]);
assign l_36[100]    = ( l_37 [100]);
assign l_36[101]    = ( l_37 [101]);
assign l_36[102]    = ( l_37 [102]);
assign l_36[103]    = ( l_37 [103]);
assign l_36[104]    = ( l_37 [104]);
assign l_36[105]    = ( l_37 [105]);
assign l_36[106]    = ( l_37 [106]);
assign l_36[107]    = ( l_37 [107]);
assign l_36[108]    = ( l_37 [108]);
assign l_36[109]    = ( l_37 [109]);
assign l_36[110]    = ( l_37 [110]);
assign l_36[111]    = ( l_37 [111]);
assign l_36[112]    = ( l_37 [112]);
assign l_36[113]    = ( l_37 [113]);
assign l_36[114]    = ( l_37 [114]);
assign l_36[115]    = ( l_37 [115]);
assign l_36[116]    = ( l_37 [116]);
assign l_36[117]    = ( l_37 [117]);
assign l_36[118]    = ( l_37 [118]);
assign l_36[119]    = ( l_37 [119]);
assign l_36[120]    = ( l_37 [120]);
assign l_36[121]    = ( l_37 [121]);
assign l_36[122]    = ( l_37 [122]);
assign l_36[123]    = ( l_37 [123]);
assign l_36[124]    = ( l_37 [124]);
assign l_36[125]    = ( l_37 [125]);
assign l_36[126]    = ( l_37 [126]);
assign l_36[127]    = ( l_37 [127]);
assign l_36[128]    = ( l_37 [128]);
assign l_36[129]    = ( l_37 [129]);
assign l_36[130]    = ( l_37 [130]);
assign l_36[131]    = ( l_37 [131]);
assign l_36[132]    = ( l_37 [132]);
assign l_36[133]    = ( l_37 [133]);
assign l_36[134]    = ( l_37 [134]);
assign l_36[135]    = ( l_37 [135]);
assign l_36[136]    = ( l_37 [136]);
assign l_36[137]    = ( l_37 [137]);
assign l_36[138]    = ( l_37 [138]);
assign l_36[139]    = ( l_37 [139]);
assign l_36[140]    = ( l_37 [140]);
assign l_36[141]    = ( l_37 [141]);
assign l_36[142]    = ( l_37 [142]);
assign l_36[143]    = ( l_37 [143]);
assign l_36[144]    = ( l_37 [144]);
assign l_36[145]    = ( l_37 [145]);
assign l_36[146]    = ( l_37 [146]);
assign l_36[147]    = ( l_37 [147]);
assign l_36[148]    = ( l_37 [148]);
assign l_36[149]    = ( l_37 [149]);
assign l_36[150]    = ( l_37 [150]);
assign l_36[151]    = ( l_37 [151]);
assign l_36[152]    = ( l_37 [152]);
assign l_36[153]    = ( l_37 [153]);
assign l_36[154]    = ( l_37 [154]);
assign l_36[155]    = ( l_37 [155]);
assign l_36[156]    = ( l_37 [156]);
assign l_36[157]    = ( l_37 [157]);
assign l_36[158]    = ( l_37 [158]);
assign l_36[159]    = ( l_37 [159]);
assign l_36[160]    = ( l_37 [160]);
assign l_36[161]    = ( l_37 [161]);
assign l_36[162]    = ( l_37 [162]);
assign l_36[163]    = ( l_37 [163]);
assign l_36[164]    = ( l_37 [164]);
assign l_36[165]    = ( l_37 [165]);
assign l_36[166]    = ( l_37 [166]);
assign l_36[167]    = ( l_37 [167]);
assign l_36[168]    = ( l_37 [168]);
assign l_36[169]    = ( l_37 [169]);
assign l_36[170]    = ( l_37 [170]);
assign l_36[171]    = ( l_37 [171]);
assign l_36[172]    = ( l_37 [172]);
assign l_36[173]    = ( l_37 [173]);
assign l_36[174]    = ( l_37 [174]);
assign l_36[175]    = ( l_37 [175]);
assign l_36[176]    = ( l_37 [176]);
assign l_36[177]    = ( l_37 [177]);
assign l_36[178]    = ( l_37 [178]);
assign l_36[179]    = ( l_37 [179]);
assign l_36[180]    = ( l_37 [180]);
assign l_36[181]    = ( l_37 [181]);
assign l_36[182]    = ( l_37 [182]);
assign l_36[183]    = ( l_37 [183]);
assign l_36[184]    = ( l_37 [184]);
assign l_36[185]    = ( l_37 [185]);
assign l_36[186]    = ( l_37 [186]);
assign l_36[187]    = ( l_37 [187]);
assign l_36[188]    = ( l_37 [188]);
assign l_36[189]    = ( l_37 [189]);
assign l_36[190]    = ( l_37 [190]);
assign l_36[191]    = ( l_37 [191]);
assign l_36[192]    = ( l_37 [192]);
assign l_36[193]    = ( l_37 [193]);
assign l_36[194]    = ( l_37 [194]);
assign l_36[195]    = ( l_37 [195]);
assign l_36[196]    = ( l_37 [196]);
assign l_36[197]    = ( l_37 [197]);
assign l_36[198]    = ( l_37 [198]);
assign l_36[199]    = ( l_37 [199]);
assign l_36[200]    = ( l_37 [200]);
assign l_36[201]    = ( l_37 [201]);
assign l_36[202]    = ( l_37 [202]);
assign l_36[203]    = ( l_37 [203]);
assign l_36[204]    = ( l_37 [204]);
assign l_36[205]    = ( l_37 [205]);
assign l_36[206]    = ( l_37 [206]);
assign l_36[207]    = ( l_37 [207]);
assign l_36[208]    = ( l_37 [208]);
assign l_36[209]    = ( l_37 [209]);
assign l_36[210]    = ( l_37 [210]);
assign l_36[211]    = ( l_37 [211]);
assign l_36[212]    = ( l_37 [212]);
assign l_36[213]    = ( l_37 [213]);
assign l_36[214]    = ( l_37 [214]);
assign l_36[215]    = ( l_37 [215]);
assign l_36[216]    = ( l_37 [216]);
assign l_36[217]    = ( l_37 [217]);
assign l_36[218]    = ( l_37 [218]);
assign l_36[219]    = ( l_37 [219]);
assign l_36[220]    = ( l_37 [220]);
assign l_36[221]    = ( l_37 [221]);
assign l_36[222]    = ( l_37 [222]);
assign l_36[223]    = ( l_37 [223]);
assign l_36[224]    = ( l_37 [224]);
assign l_36[225]    = ( l_37 [225]);
assign l_36[226]    = ( l_37 [226]);
assign l_36[227]    = ( l_37 [227]);
assign l_36[228]    = ( l_37 [228]);
assign l_36[229]    = ( l_37 [229]);
assign l_36[230]    = ( l_37 [230]);
assign l_36[231]    = ( l_37 [231]);
assign l_36[232]    = ( l_37 [232]);
assign l_36[233]    = ( l_37 [233]);
assign l_36[234]    = ( l_37 [234]);
assign l_36[235]    = ( l_37 [235]);
assign l_36[236]    = ( l_37 [236]);
assign l_36[237]    = ( l_37 [237]);
assign l_36[238]    = ( l_37 [238]);
assign l_36[239]    = ( l_37 [239]);
assign l_36[240]    = ( l_37 [240]);
assign l_36[241]    = ( l_37 [241]);
assign l_36[242]    = ( l_37 [242]);
assign l_36[243]    = ( l_37 [243]);
assign l_36[244]    = ( l_37 [244]);
assign l_36[245]    = ( l_37 [245]);
assign l_36[246]    = ( l_37 [246]);
assign l_36[247]    = ( l_37 [247]);
assign l_36[248]    = ( l_37 [248]);
assign l_36[249]    = ( l_37 [249]);
assign l_36[250]    = ( l_37 [250]);
assign l_36[251]    = ( l_37 [251]);
assign l_36[252]    = ( l_37 [252]);
assign l_36[253]    = ( l_37 [253]);
assign l_36[254]    = ( l_37 [254]);
assign l_36[255]    = ( l_37 [255]);
assign l_36[256]    = ( l_37 [256]);
assign l_36[257]    = ( l_37 [257]);
assign l_36[258]    = ( l_37 [258]);
assign l_36[259]    = ( l_37 [259]);
assign l_36[260]    = ( l_37 [260]);
assign l_36[261]    = ( l_37 [261]);
assign l_36[262]    = ( l_37 [262]);
assign l_36[263]    = ( l_37 [263]);
assign l_36[264]    = ( l_37 [264]);
assign l_36[265]    = ( l_37 [265]);
assign l_36[266]    = ( l_37 [266]);
assign l_36[267]    = ( l_37 [267]);
assign l_36[268]    = ( l_37 [268]);
assign l_36[269]    = ( l_37 [269]);
assign l_36[270]    = ( l_37 [270]);
assign l_36[271]    = ( l_37 [271]);
assign l_36[272]    = ( l_37 [272]);
assign l_36[273]    = ( l_37 [273]);
assign l_36[274]    = ( l_37 [274]);
assign l_36[275]    = ( l_37 [275]);
assign l_36[276]    = ( l_37 [276]);
assign l_36[277]    = ( l_37 [277]);
assign l_36[278]    = ( l_37 [278]);
assign l_36[279]    = ( l_37 [279]);
assign l_36[280]    = ( l_37 [280]);
assign l_36[281]    = ( l_37 [281]);
assign l_36[282]    = ( l_37 [282]);
assign l_36[283]    = ( l_37 [283]);
assign l_36[284]    = ( l_37 [284]);
assign l_36[285]    = ( l_37 [285]);
assign l_36[286]    = ( l_37 [286]);
assign l_36[287]    = ( l_37 [287]);
assign l_36[288]    = ( l_37 [288]);
assign l_36[289]    = ( l_37 [289]);
assign l_36[290]    = ( l_37 [290]);
assign l_36[291]    = ( l_37 [291]);
assign l_36[292]    = ( l_37 [292]);
assign l_36[293]    = ( l_37 [293]);
assign l_36[294]    = ( l_37 [294]);
assign l_36[295]    = ( l_37 [295]);
assign l_36[296]    = ( l_37 [296]);
assign l_36[297]    = ( l_37 [297]);
assign l_36[298]    = ( l_37 [298]);
assign l_36[299]    = ( l_37 [299]);
assign l_36[300]    = ( l_37 [300]);
assign l_36[301]    = ( l_37 [301]);
assign l_36[302]    = ( l_37 [302]);
assign l_36[303]    = ( l_37 [303]);
assign l_36[304]    = ( l_37 [304]);
assign l_36[305]    = ( l_37 [305]);
assign l_36[306]    = ( l_37 [306]);
assign l_36[307]    = ( l_37 [307]);
assign l_36[308]    = ( l_37 [308]);
assign l_36[309]    = ( l_37 [309]);
assign l_36[310]    = ( l_37 [310]);
assign l_36[311]    = ( l_37 [311]);
assign l_36[312]    = ( l_37 [312]);
assign l_36[313]    = ( l_37 [313]);
assign l_36[314]    = ( l_37 [314]);
assign l_36[315]    = ( l_37 [315]);
assign l_36[316]    = ( l_37 [316]);
assign l_36[317]    = ( l_37 [317]);
assign l_36[318]    = ( l_37 [318]);
assign l_36[319]    = ( l_37 [319]);
assign l_36[320]    = ( l_37 [320]);
assign l_36[321]    = ( l_37 [321]);
assign l_36[322]    = ( l_37 [322]);
assign l_36[323]    = ( l_37 [323]);
assign l_36[324]    = ( l_37 [324]);
assign l_36[325]    = ( l_37 [325]);
assign l_36[326]    = ( l_37 [326]);
assign l_36[327]    = ( l_37 [327]);
assign l_36[328]    = ( l_37 [328]);
assign l_36[329]    = ( l_37 [329]);
assign l_36[330]    = ( l_37 [330]);
assign l_36[331]    = ( l_37 [331]);
assign l_36[332]    = ( l_37 [332]);
assign l_36[333]    = ( l_37 [333]);
assign l_36[334]    = ( l_37 [334]);
assign l_36[335]    = ( l_37 [335]);
assign l_36[336]    = ( l_37 [336]);
assign l_36[337]    = ( l_37 [337]);
assign l_36[338]    = ( l_37 [338]);
assign l_36[339]    = ( l_37 [339]);
assign l_36[340]    = ( l_37 [340]);
assign l_36[341]    = ( l_37 [341]);
assign l_36[342]    = ( l_37 [342]);
assign l_36[343]    = ( l_37 [343]);
assign l_36[344]    = ( l_37 [344]);
assign l_36[345]    = ( l_37 [345]);
assign l_36[346]    = ( l_37 [346]);
assign l_36[347]    = ( l_37 [347]);
assign l_36[348]    = ( l_37 [348]);
assign l_36[349]    = ( l_37 [349]);
assign l_36[350]    = ( l_37 [350]);
assign l_36[351]    = ( l_37 [351]);
assign l_36[352]    = ( l_37 [352]);
assign l_36[353]    = ( l_37 [353]);
assign l_36[354]    = ( l_37 [354]);
assign l_36[355]    = ( l_37 [355]);
assign l_36[356]    = ( l_37 [356]);
assign l_36[357]    = ( l_37 [357]);
assign l_36[358]    = ( l_37 [358]);
assign l_36[359]    = ( l_37 [359]);
assign l_36[360]    = ( l_37 [360]);
assign l_36[361]    = ( l_37 [361]);
assign l_36[362]    = ( l_37 [362]);
assign l_36[363]    = ( l_37 [363]);
assign l_36[364]    = ( l_37 [364]);
assign l_36[365]    = ( l_37 [365]);
assign l_36[366]    = ( l_37 [366]);
assign l_36[367]    = ( l_37 [367]);
assign l_36[368]    = ( l_37 [368]);
assign l_36[369]    = ( l_37 [369]);
assign l_36[370]    = ( l_37 [370]);
assign l_36[371]    = ( l_37 [371]);
assign l_36[372]    = ( l_37 [372]);
assign l_36[373]    = ( l_37 [373]);
assign l_36[374]    = ( l_37 [374]);
assign l_36[375]    = ( l_37 [375]);
assign l_36[376]    = ( l_37 [376]);
assign l_36[377]    = ( l_37 [377]);
assign l_36[378]    = ( l_37 [378]);
assign l_36[379]    = ( l_37 [379]);
assign l_36[380]    = ( l_37 [380]);
assign l_36[381]    = ( l_37 [381]);
assign l_36[382]    = ( l_37 [382]);
assign l_36[383]    = ( l_37 [383]);
assign l_36[384]    = ( l_37 [384]);
assign l_36[385]    = ( l_37 [385]);
assign l_36[386]    = ( l_37 [386]);
assign l_36[387]    = ( l_37 [387]);
assign l_36[388]    = ( l_37 [388]);
assign l_36[389]    = ( l_37 [389]);
assign l_36[390]    = ( l_37 [390]);
assign l_36[391]    = ( l_37 [391]);
assign l_36[392]    = ( l_37 [392]);
assign l_36[393]    = ( l_37 [393]);
assign l_36[394]    = ( l_37 [394]);
assign l_36[395]    = ( l_37 [395]);
assign l_36[396]    = ( l_37 [396]);
assign l_36[397]    = ( l_37 [397]);
assign l_36[398]    = ( l_37 [398]);
assign l_36[399]    = ( l_37 [399]);
assign l_36[400]    = ( l_37 [400]);
assign l_36[401]    = ( l_37 [401]);
assign l_36[402]    = ( l_37 [402]);
assign l_36[403]    = ( l_37 [403]);
assign l_36[404]    = ( l_37 [404]);
assign l_36[405]    = ( l_37 [405]);
assign l_36[406]    = ( l_37 [406]);
assign l_36[407]    = ( l_37 [407]);
assign l_36[408]    = ( l_37 [408]);
assign l_36[409]    = ( l_37 [409]);
assign l_36[410]    = ( l_37 [410]);
assign l_36[411]    = ( l_37 [411]);
assign l_36[412]    = ( l_37 [412]);
assign l_36[413]    = ( l_37 [413]);
assign l_36[414]    = ( l_37 [414]);
assign l_36[415]    = ( l_37 [415]);
assign l_36[416]    = ( l_37 [416]);
assign l_36[417]    = ( l_37 [417]);
assign l_36[418]    = ( l_37 [418]);
assign l_36[419]    = ( l_37 [419]);
assign l_36[420]    = ( l_37 [420]);
assign l_36[421]    = ( l_37 [421]);
assign l_36[422]    = ( l_37 [422]);
assign l_36[423]    = ( l_37 [423]);
assign l_36[424]    = ( l_37 [424]);
assign l_36[425]    = ( l_37 [425]);
assign l_36[426]    = ( l_37 [426]);
assign l_36[427]    = ( l_37 [427]);
assign l_36[428]    = ( l_37 [428]);
assign l_36[429]    = ( l_37 [429]);
assign l_36[430]    = ( l_37 [430]);
assign l_36[431]    = ( l_37 [431]);
assign l_36[432]    = ( l_37 [432]);
assign l_36[433]    = ( l_37 [433]);
assign l_36[434]    = ( l_37 [434]);
assign l_36[435]    = ( l_37 [435]);
assign l_36[436]    = ( l_37 [436]);
assign l_36[437]    = ( l_37 [437]);
assign l_36[438]    = ( l_37 [438]);
assign l_36[439]    = ( l_37 [439]);
assign l_36[440]    = ( l_37 [440]);
assign l_36[441]    = ( l_37 [441]);
assign l_36[442]    = ( l_37 [442]);
assign l_36[443]    = ( l_37 [443]);
assign l_36[444]    = ( l_37 [444]);
assign l_36[445]    = ( l_37 [445]);
assign l_36[446]    = ( l_37 [446]);
assign l_36[447]    = ( l_37 [447]);
assign l_36[448]    = ( l_37 [448]);
assign l_36[449]    = ( l_37 [449]);
assign l_36[450]    = ( l_37 [450]);
assign l_36[451]    = ( l_37 [451]);
assign l_36[452]    = ( l_37 [452]);
assign l_36[453]    = ( l_37 [453]);
assign l_36[454]    = ( l_37 [454]);
assign l_36[455]    = ( l_37 [455]);
assign l_36[456]    = ( l_37 [456]);
assign l_36[457]    = ( l_37 [457]);
assign l_36[458]    = ( l_37 [458]);
assign l_36[459]    = ( l_37 [459]);
assign l_36[460]    = ( l_37 [460]);
assign l_36[461]    = ( l_37 [461]);
assign l_36[462]    = ( l_37 [462]);
assign l_36[463]    = ( l_37 [463]);
assign l_36[464]    = ( l_37 [464]);
assign l_36[465]    = ( l_37 [465]);
assign l_36[466]    = ( l_37 [466]);
assign l_36[467]    = ( l_37 [467]);
assign l_36[468]    = ( l_37 [468]);
assign l_36[469]    = ( l_37 [469]);
assign l_36[470]    = ( l_37 [470]);
assign l_36[471]    = ( l_37 [471]);
assign l_36[472]    = ( l_37 [472]);
assign l_36[473]    = ( l_37 [473]);
assign l_36[474]    = ( l_37 [474]);
assign l_36[475]    = ( l_37 [475]);
assign l_36[476]    = ( l_37 [476]);
assign l_36[477]    = ( l_37 [477]);
assign l_36[478]    = ( l_37 [478]);
assign l_36[479]    = ( l_37 [479]);
assign l_36[480]    = ( l_37 [480]);
assign l_36[481]    = ( l_37 [481]);
assign l_36[482]    = ( l_37 [482]);
assign l_36[483]    = ( l_37 [483]);
assign l_36[484]    = ( l_37 [484]);
assign l_36[485]    = ( l_37 [485]);
assign l_36[486]    = ( l_37 [486]);
assign l_36[487]    = ( l_37 [487]);
assign l_36[488]    = ( l_37 [488]);
assign l_36[489]    = ( l_37 [489]);
assign l_36[490]    = ( l_37 [490]);
assign l_36[491]    = ( l_37 [491]);
assign l_36[492]    = ( l_37 [492]);
assign l_36[493]    = ( l_37 [493]);
assign l_36[494]    = ( l_37 [494]);
assign l_36[495]    = ( l_37 [495]);
assign l_36[496]    = ( l_37 [496]);
assign l_36[497]    = ( l_37 [497]);
assign l_36[498]    = ( l_37 [498]);
assign l_36[499]    = ( l_37 [499]);
assign l_36[500]    = ( l_37 [500]);
assign l_36[501]    = ( l_37 [501]);
assign l_36[502]    = ( l_37 [502]);
assign l_36[503]    = ( l_37 [503]);
assign l_36[504]    = ( l_37 [504]);
assign l_36[505]    = ( l_37 [505]);
assign l_36[506]    = ( l_37 [506]);
assign l_36[507]    = ( l_37 [507]);
assign l_36[508]    = ( l_37 [508]);
assign l_36[509]    = ( l_37 [509]);
assign l_36[510]    = ( l_37 [510]);
assign l_36[511]    = ( l_37 [511]);
assign l_36[512]    = ( l_37 [512]);
assign l_36[513]    = ( l_37 [513]);
assign l_36[514]    = ( l_37 [514]);
assign l_36[515]    = ( l_37 [515]);
assign l_36[516]    = ( l_37 [516]);
assign l_36[517]    = ( l_37 [517]);
assign l_36[518]    = ( l_37 [518]);
assign l_36[519]    = ( l_37 [519]);
assign l_36[520]    = ( l_37 [520]);
assign l_36[521]    = ( l_37 [521]);
assign l_36[522]    = ( l_37 [522]);
assign l_36[523]    = ( l_37 [523]);
assign l_36[524]    = ( l_37 [524]);
assign l_36[525]    = ( l_37 [525]);
assign l_36[526]    = ( l_37 [526]);
assign l_36[527]    = ( l_37 [527]);
assign l_36[528]    = ( l_37 [528]);
assign l_36[529]    = ( l_37 [529]);
assign l_36[530]    = ( l_37 [530] & !i[1800]) | ( l_37 [531] &  i[1800]);
assign l_36[531]    = ( l_37 [532] & !i[1800]) | ( l_37 [533] &  i[1800]);
assign l_36[532]    = ( l_37 [534] & !i[1800]) | ( l_37 [535] &  i[1800]);
assign l_36[533]    = ( l_37 [536] & !i[1800]) | ( l_37 [537] &  i[1800]);
assign l_36[534]    = ( l_37 [538] & !i[1800]) | ( l_37 [539] &  i[1800]);
assign l_36[535]    = ( l_37 [540] & !i[1800]) | ( l_37 [541] &  i[1800]);
assign l_36[536]    = ( l_37 [542] & !i[1800]) | ( l_37 [543] &  i[1800]);
assign l_36[537]    = ( l_37 [544] & !i[1800]) | ( l_37 [545] &  i[1800]);
assign l_36[538]    = ( l_37 [546] & !i[1800]) | ( l_37 [547] &  i[1800]);
assign l_36[539]    = ( l_37 [548] & !i[1800]) | ( l_37 [549] &  i[1800]);
assign l_36[540]    = ( l_37 [550] & !i[1800]) | ( l_37 [551] &  i[1800]);
assign l_36[541]    = ( l_37 [552] & !i[1800]) | ( l_37 [553] &  i[1800]);
assign l_36[542]    = ( l_37 [554] & !i[1800]) | ( l_37 [555] &  i[1800]);
assign l_36[543]    = ( l_37 [556] & !i[1800]) | ( l_37 [557] &  i[1800]);
assign l_36[544]    = ( l_37 [558] & !i[1800]) | ( l_37 [559] &  i[1800]);
assign l_36[545]    = ( l_37 [560] & !i[1800]) | ( l_37 [561] &  i[1800]);
assign l_36[546]    = ( l_37 [562] & !i[1800]) | ( l_37 [563] &  i[1800]);
assign l_36[547]    = ( l_37 [564] & !i[1800]) | ( l_37 [565] &  i[1800]);
assign l_36[548]    = ( l_37 [566] & !i[1800]) | ( l_37 [567] &  i[1800]);
assign l_36[549]    = ( l_37 [568] & !i[1800]) | ( l_37 [569] &  i[1800]);
assign l_36[550]    = ( l_37 [570] & !i[1800]) | ( l_37 [571] &  i[1800]);
assign l_36[551]    = ( l_37 [572] & !i[1800]) | ( l_37 [573] &  i[1800]);
assign l_36[552]    = ( l_37 [574] & !i[1800]) | ( l_37 [575] &  i[1800]);
assign l_36[553]    = ( l_37 [576] & !i[1800]) | ( l_37 [577] &  i[1800]);
assign l_36[554]    = ( l_37 [578] & !i[1800]) | ( l_37 [579] &  i[1800]);
assign l_36[555]    = ( l_37 [580] & !i[1800]) | ( l_37 [581] &  i[1800]);
assign l_36[556]    = ( l_37 [582] & !i[1800]) | ( l_37 [583] &  i[1800]);
assign l_36[557]    = ( l_37 [584] & !i[1800]) | ( l_37 [585] &  i[1800]);
assign l_36[558]    = ( l_37 [586] & !i[1800]) | ( l_37 [587] &  i[1800]);
assign l_36[559]    = ( l_37 [588] & !i[1800]) | ( l_37 [589] &  i[1800]);
assign l_36[560]    = ( l_37 [590] & !i[1800]) | ( l_37 [591] &  i[1800]);
assign l_36[561]    = ( l_37 [592] & !i[1800]) | ( l_37 [593] &  i[1800]);
assign l_36[562]    = ( l_37 [594] & !i[1800]) | ( l_37 [595] &  i[1800]);
assign l_36[563]    = ( l_37 [596] & !i[1800]) | ( l_37 [597] &  i[1800]);
assign l_36[564]    = ( l_37 [598] & !i[1800]) | ( l_37 [599] &  i[1800]);
assign l_36[565]    = ( l_37 [600] & !i[1800]) | ( l_37 [601] &  i[1800]);
assign l_36[566]    = ( l_37 [602] & !i[1800]) | ( l_37 [603] &  i[1800]);
assign l_36[567]    = ( l_37 [604] & !i[1800]) | ( l_37 [605] &  i[1800]);
assign l_36[568]    = ( l_37 [606] & !i[1800]) | ( l_37 [607] &  i[1800]);
assign l_36[569]    = ( l_37 [608] & !i[1800]) | ( l_37 [609] &  i[1800]);
assign l_36[570]    = ( l_37 [610] & !i[1800]) | ( l_37 [611] &  i[1800]);
assign l_36[571]    = ( l_37 [612] & !i[1800]) | ( l_37 [613] &  i[1800]);
assign l_36[572]    = ( l_37 [614] & !i[1800]) | ( l_37 [615] &  i[1800]);
assign l_36[573]    = ( l_37 [616] & !i[1800]) | ( l_37 [617] &  i[1800]);
assign l_36[574]    = ( l_37 [618] & !i[1800]) | ( l_37 [619] &  i[1800]);
assign l_36[575]    = ( l_37 [620] & !i[1800]) | ( l_37 [621] &  i[1800]);
assign l_36[576]    = ( l_37 [622] & !i[1800]) | ( l_37 [623] &  i[1800]);
assign l_36[577]    = ( l_37 [624] & !i[1800]) | ( l_37 [625] &  i[1800]);
assign l_36[578]    = ( l_37 [626] & !i[1800]) | ( l_37 [627] &  i[1800]);
assign l_36[579]    = ( l_37 [628] & !i[1800]) | ( l_37 [629] &  i[1800]);
assign l_36[580]    = ( l_37 [630] & !i[1800]) | ( l_37 [631] &  i[1800]);
assign l_36[581]    = ( l_37 [632] & !i[1800]) | ( l_37 [633] &  i[1800]);
assign l_36[582]    = ( l_37 [634] & !i[1800]) | ( l_37 [635] &  i[1800]);
assign l_36[583]    = ( l_37 [636] & !i[1800]) | ( l_37 [637] &  i[1800]);
assign l_36[584]    = ( l_37 [638] & !i[1800]) | ( l_37 [639] &  i[1800]);
assign l_36[585]    = ( l_37 [640] & !i[1800]) | ( l_37 [641] &  i[1800]);
assign l_36[586]    = ( l_37 [642] & !i[1800]) | ( l_37 [643] &  i[1800]);
assign l_36[587]    = ( l_37 [644] & !i[1800]) | ( l_37 [645] &  i[1800]);
assign l_36[588]    = ( l_37 [646] & !i[1800]) | ( l_37 [647] &  i[1800]);
assign l_36[589]    = ( l_37 [648] & !i[1800]) | ( l_37 [649] &  i[1800]);
assign l_36[590]    = ( l_37 [650] & !i[1800]) | ( l_37 [651] &  i[1800]);
assign l_36[591]    = ( l_37 [652] & !i[1800]) | ( l_37 [653] &  i[1800]);
assign l_36[592]    = ( l_37 [654] & !i[1800]) | ( l_37 [655] &  i[1800]);
assign l_36[593]    = ( l_37 [656] & !i[1800]) | ( l_37 [657] &  i[1800]);
assign l_36[594]    = ( l_37 [658] & !i[1800]) | ( l_37 [659] &  i[1800]);
assign l_36[595]    = ( l_37 [660] & !i[1800]) | ( l_37 [661] &  i[1800]);
assign l_36[596]    = ( l_37 [662] & !i[1800]) | ( l_37 [663] &  i[1800]);
assign l_36[597]    = ( l_37 [664] & !i[1800]) | ( l_37 [665] &  i[1800]);
assign l_36[598]    = ( l_37 [666] & !i[1800]) | ( l_37 [667] &  i[1800]);
assign l_36[599]    = ( l_37 [668] & !i[1800]) | ( l_37 [669] &  i[1800]);
assign l_36[600]    = ( l_37 [670] & !i[1800]) | ( l_37 [671] &  i[1800]);
assign l_36[601]    = ( l_37 [672] & !i[1800]) | ( l_37 [673] &  i[1800]);
assign l_36[602]    = ( l_37 [674] & !i[1800]) | ( l_37 [675] &  i[1800]);
assign l_36[603]    = ( l_37 [676] & !i[1800]) | ( l_37 [677] &  i[1800]);
assign l_36[604]    = ( l_37 [678] & !i[1800]) | ( l_37 [679] &  i[1800]);
assign l_36[605]    = ( l_37 [680] & !i[1800]) | ( l_37 [681] &  i[1800]);
assign l_36[606]    = ( l_37 [682] & !i[1800]) | ( l_37 [683] &  i[1800]);
assign l_36[607]    = ( l_37 [684] & !i[1800]) | ( l_37 [685] &  i[1800]);
assign l_36[608]    = ( l_37 [686] & !i[1800]) | ( l_37 [687] &  i[1800]);
assign l_36[609]    = ( l_37 [688] & !i[1800]) | ( l_37 [689] &  i[1800]);
assign l_36[610]    = ( l_37 [690] & !i[1800]) | ( l_37 [691] &  i[1800]);
assign l_36[611]    = ( l_37 [692] & !i[1800]) | ( l_37 [693] &  i[1800]);
assign l_36[612]    = ( l_37 [694] & !i[1800]) | ( l_37 [695] &  i[1800]);
assign l_36[613]    = ( l_37 [696] & !i[1800]) | ( l_37 [697] &  i[1800]);
assign l_36[614]    = ( l_37 [698] & !i[1800]) | ( l_37 [699] &  i[1800]);
assign l_36[615]    = ( l_37 [700] & !i[1800]) | ( l_37 [701] &  i[1800]);
assign l_36[616]    = ( l_37 [702] & !i[1800]) | ( l_37 [703] &  i[1800]);
assign l_36[617]    = ( l_37 [704] & !i[1800]) | ( l_37 [705] &  i[1800]);
assign l_36[618]    = ( l_37 [706] & !i[1800]) | ( l_37 [707] &  i[1800]);
assign l_36[619]    = ( l_37 [708] & !i[1800]) | ( l_37 [709] &  i[1800]);
assign l_36[620]    = ( l_37 [710] & !i[1800]) | ( l_37 [711] &  i[1800]);
assign l_36[621]    = ( l_37 [712] & !i[1800]) | ( l_37 [713] &  i[1800]);
assign l_36[622]    = ( l_37 [714] & !i[1800]) | ( l_37 [715] &  i[1800]);
assign l_36[623]    = ( l_37 [716] & !i[1800]) | ( l_37 [717] &  i[1800]);
assign l_36[624]    = ( l_37 [718] & !i[1800]) | ( l_37 [719] &  i[1800]);
assign l_36[625]    = ( l_37 [720] & !i[1800]) | ( l_37 [721] &  i[1800]);
assign l_36[626]    = ( l_37 [722] & !i[1800]) | ( l_37 [723] &  i[1800]);
assign l_36[627]    = ( l_37 [724] & !i[1800]) | ( l_37 [725] &  i[1800]);
assign l_36[628]    = ( l_37 [726] & !i[1800]) | ( l_37 [727] &  i[1800]);
assign l_36[629]    = ( l_37 [728] & !i[1800]) | ( l_37 [729] &  i[1800]);
assign l_36[630]    = ( l_37 [730] & !i[1800]) | ( l_37 [731] &  i[1800]);
assign l_36[631]    = ( l_37 [732] & !i[1800]) | ( l_37 [733] &  i[1800]);
assign l_36[632]    = ( l_37 [734] & !i[1800]) | ( l_37 [735] &  i[1800]);
assign l_36[633]    = ( l_37 [736] & !i[1800]) | ( l_37 [737] &  i[1800]);
assign l_36[634]    = ( l_37 [738] & !i[1800]) | ( l_37 [739] &  i[1800]);
assign l_36[635]    = ( l_37 [740] & !i[1800]) | ( l_37 [741] &  i[1800]);
assign l_36[636]    = ( l_37 [742] & !i[1800]) | ( l_37 [743] &  i[1800]);
assign l_36[637]    = ( l_37 [744] & !i[1800]) | ( l_37 [745] &  i[1800]);
assign l_36[638]    = ( l_37 [746] & !i[1800]) | ( l_37 [747] &  i[1800]);
assign l_36[639]    = ( l_37 [748] & !i[1800]) | ( l_37 [749] &  i[1800]);
assign l_36[640]    = ( l_37 [750] & !i[1800]) | ( l_37 [751] &  i[1800]);
assign l_36[641]    = ( l_37 [752] & !i[1800]) | ( l_37 [753] &  i[1800]);
assign l_36[642]    = ( l_37 [754] & !i[1800]) | ( l_37 [755] &  i[1800]);
assign l_36[643]    = ( l_37 [756] & !i[1800]) | ( l_37 [757] &  i[1800]);
assign l_36[644]    = ( l_37 [758] & !i[1800]) | ( l_37 [759] &  i[1800]);
assign l_36[645]    = ( l_37 [760] & !i[1800]) | ( l_37 [761] &  i[1800]);
assign l_36[646]    = ( l_37 [762] & !i[1800]) | ( l_37 [763] &  i[1800]);
assign l_36[647]    = ( l_37 [764] & !i[1800]) | ( l_37 [765] &  i[1800]);
assign l_36[648]    = ( l_37 [766] & !i[1800]) | ( l_37 [767] &  i[1800]);
assign l_36[649]    = ( l_37 [768] & !i[1800]) | ( l_37 [769] &  i[1800]);
assign l_36[650]    = ( l_37 [770] & !i[1800]) | ( l_37 [771] &  i[1800]);
assign l_36[651]    = ( l_37 [772] & !i[1800]) | ( l_37 [773] &  i[1800]);
assign l_36[652]    = ( l_37 [774] & !i[1800]) | ( l_37 [775] &  i[1800]);
assign l_36[653]    = ( l_37 [776] & !i[1800]) | ( l_37 [777] &  i[1800]);
assign l_36[654]    = ( l_37 [778] & !i[1800]) | ( l_37 [779] &  i[1800]);
assign l_36[655]    = ( l_37 [780] & !i[1800]) | ( l_37 [781] &  i[1800]);
assign l_36[656]    = ( l_37 [782] & !i[1800]) | ( l_37 [783] &  i[1800]);
assign l_36[657]    = ( l_37 [784] & !i[1800]) | ( l_37 [785] &  i[1800]);
assign l_36[658]    = ( l_37 [786] & !i[1800]) | ( l_37 [787] &  i[1800]);
assign l_36[659]    = ( l_37 [788] & !i[1800]) | ( l_37 [789] &  i[1800]);
assign l_36[660]    = ( l_37 [790] & !i[1800]) | ( l_37 [791] &  i[1800]);
assign l_36[661]    = ( l_37 [792] & !i[1800]) | ( l_37 [793] &  i[1800]);
assign l_36[662]    = ( l_37 [794] & !i[1800]) | ( l_37 [795] &  i[1800]);
assign l_36[663]    = ( l_37 [796] & !i[1800]) | ( l_37 [797] &  i[1800]);
assign l_36[664]    = ( l_37 [798] & !i[1800]) | ( l_37 [799] &  i[1800]);
assign l_36[665]    = ( l_37 [800] & !i[1800]) | ( l_37 [801] &  i[1800]);
assign l_36[666]    = ( l_37 [802] & !i[1800]) | ( l_37 [803] &  i[1800]);
assign l_36[667]    = ( l_37 [804] & !i[1800]) | ( l_37 [805] &  i[1800]);
assign l_36[668]    = ( l_37 [806] & !i[1800]) | ( l_37 [807] &  i[1800]);
assign l_36[669]    = ( l_37 [808] & !i[1800]) | ( l_37 [809] &  i[1800]);
assign l_36[670]    = ( l_37 [810] & !i[1800]) | ( l_37 [811] &  i[1800]);
assign l_36[671]    = ( l_37 [812] & !i[1800]) | ( l_37 [813] &  i[1800]);
assign l_36[672]    = ( l_37 [814] & !i[1800]) | ( l_37 [815] &  i[1800]);
assign l_36[673]    = ( l_37 [816] & !i[1800]) | ( l_37 [817] &  i[1800]);
assign l_36[674]    = ( l_37 [818] & !i[1800]) | ( l_37 [819] &  i[1800]);
assign l_36[675]    = ( l_37 [820] & !i[1800]) | ( l_37 [821] &  i[1800]);
assign l_36[676]    = ( l_37 [822] & !i[1800]) | ( l_37 [823] &  i[1800]);
assign l_36[677]    = ( l_37 [824] & !i[1800]) | ( l_37 [825] &  i[1800]);
assign l_36[678]    = ( l_37 [826] & !i[1800]) | ( l_37 [827] &  i[1800]);
assign l_36[679]    = ( l_37 [828] & !i[1800]) | ( l_37 [829] &  i[1800]);
assign l_36[680]    = ( l_37 [830] & !i[1800]) | ( l_37 [831] &  i[1800]);
assign l_36[681]    = ( l_37 [832] & !i[1800]) | ( l_37 [833] &  i[1800]);
assign l_36[682]    = ( l_37 [834] & !i[1800]) | ( l_37 [835] &  i[1800]);
assign l_36[683]    = ( l_37 [836] & !i[1800]) | ( l_37 [837] &  i[1800]);
assign l_36[684]    = ( l_37 [838] & !i[1800]) | ( l_37 [839] &  i[1800]);
assign l_36[685]    = ( l_37 [840] & !i[1800]) | ( l_37 [841] &  i[1800]);
assign l_36[686]    = ( l_37 [842] & !i[1800]) | ( l_37 [843] &  i[1800]);
assign l_36[687]    = ( l_37 [844] & !i[1800]) | ( l_37 [845] &  i[1800]);
assign l_36[688]    = ( l_37 [846] & !i[1800]) | ( l_37 [847] &  i[1800]);
assign l_36[689]    = ( l_37 [848] & !i[1800]) | ( l_37 [849] &  i[1800]);
assign l_36[690]    = ( l_37 [850] & !i[1800]) | ( l_37 [851] &  i[1800]);
assign l_36[691]    = ( l_37 [852] & !i[1800]) | ( l_37 [853] &  i[1800]);
assign l_36[692]    = ( l_37 [854] & !i[1800]) | ( l_37 [855] &  i[1800]);
assign l_36[693]    = ( l_37 [856] & !i[1800]) | ( l_37 [857] &  i[1800]);
assign l_36[694]    = ( l_37 [858] & !i[1800]) | ( l_37 [859] &  i[1800]);
assign l_36[695]    = ( l_37 [860] & !i[1800]) | ( l_37 [861] &  i[1800]);
assign l_36[696]    = ( l_37 [862] & !i[1800]) | ( l_37 [863] &  i[1800]);
assign l_36[697]    = ( l_37 [864] & !i[1800]) | ( l_37 [865] &  i[1800]);
assign l_36[698]    = ( l_37 [866] & !i[1800]) | ( l_37 [867] &  i[1800]);
assign l_36[699]    = ( l_37 [868] & !i[1800]) | ( l_37 [869] &  i[1800]);
assign l_36[700]    = ( l_37 [870] & !i[1800]) | ( l_37 [871] &  i[1800]);
assign l_36[701]    = ( l_37 [872] & !i[1800]) | ( l_37 [873] &  i[1800]);
assign l_36[702]    = ( l_37 [874] & !i[1800]) | ( l_37 [875] &  i[1800]);
assign l_36[703]    = ( l_37 [876] & !i[1800]) | ( l_37 [877] &  i[1800]);
assign l_36[704]    = ( l_37 [878] & !i[1800]) | ( l_37 [879] &  i[1800]);
assign l_36[705]    = ( l_37 [880] & !i[1800]) | ( l_37 [881] &  i[1800]);
assign l_36[706]    = ( l_37 [882] & !i[1800]) | ( l_37 [883] &  i[1800]);
assign l_36[707]    = ( l_37 [884] & !i[1800]) | ( l_37 [885] &  i[1800]);
assign l_36[708]    = ( l_37 [886] & !i[1800]) | ( l_37 [887] &  i[1800]);
assign l_36[709]    = ( l_37 [888] & !i[1800]) | ( l_37 [889] &  i[1800]);
assign l_36[710]    = ( l_37 [890] & !i[1800]) | ( l_37 [891] &  i[1800]);
assign l_36[711]    = ( l_37 [892] & !i[1800]) | ( l_37 [893] &  i[1800]);
assign l_36[712]    = ( l_37 [894] & !i[1800]) | ( l_37 [895] &  i[1800]);
assign l_36[713]    = ( l_37 [896] & !i[1800]) | ( l_37 [897] &  i[1800]);
assign l_36[714]    = ( l_37 [898] & !i[1800]) | ( l_37 [899] &  i[1800]);
assign l_36[715]    = ( l_37 [900] & !i[1800]) | ( l_37 [901] &  i[1800]);
assign l_36[716]    = ( l_37 [902] & !i[1800]) | ( l_37 [903] &  i[1800]);
assign l_36[717]    = ( l_37 [904] & !i[1800]) | ( l_37 [905] &  i[1800]);
assign l_36[718]    = ( l_37 [906] & !i[1800]) | ( l_37 [907] &  i[1800]);
assign l_36[719]    = ( l_37 [908] & !i[1800]) | ( l_37 [909] &  i[1800]);
assign l_36[720]    = ( l_37 [910] & !i[1800]) | ( l_37 [911] &  i[1800]);
assign l_36[721]    = ( l_37 [912] & !i[1800]) | ( l_37 [913] &  i[1800]);
assign l_36[722]    = ( l_37 [914] & !i[1800]) | ( l_37 [915] &  i[1800]);
assign l_36[723]    = ( l_37 [916] & !i[1800]) | ( l_37 [917] &  i[1800]);
assign l_36[724]    = ( l_37 [918] & !i[1800]) | ( l_37 [919] &  i[1800]);
assign l_36[725]    = ( l_37 [920] & !i[1800]) | ( l_37 [921] &  i[1800]);
assign l_36[726]    = ( l_37 [922] & !i[1800]) | ( l_37 [923] &  i[1800]);
assign l_36[727]    = ( l_37 [924] & !i[1800]) | ( l_37 [925] &  i[1800]);
assign l_36[728]    = ( l_37 [926] & !i[1800]) | ( l_37 [927] &  i[1800]);
assign l_36[729]    = ( l_37 [928] & !i[1800]) | ( l_37 [929] &  i[1800]);
assign l_36[730]    = ( l_37 [930] & !i[1800]) | ( l_37 [931] &  i[1800]);
assign l_36[731]    = ( l_37 [932] & !i[1800]) | ( l_37 [933] &  i[1800]);
assign l_36[732]    = ( l_37 [934] & !i[1800]) | ( l_37 [935] &  i[1800]);
assign l_36[733]    = ( l_37 [936] & !i[1800]) | ( l_37 [937] &  i[1800]);
assign l_36[734]    = ( l_37 [938] & !i[1800]) | ( l_37 [939] &  i[1800]);
assign l_36[735]    = ( l_37 [940] & !i[1800]) | ( l_37 [941] &  i[1800]);
assign l_36[736]    = ( l_37 [942] & !i[1800]) | ( l_37 [943] &  i[1800]);
assign l_36[737]    = ( l_37 [944] & !i[1800]) | ( l_37 [945] &  i[1800]);
assign l_36[738]    = ( l_37 [946] & !i[1800]) | ( l_37 [947] &  i[1800]);
assign l_36[739]    = ( l_37 [948] & !i[1800]) | ( l_37 [949] &  i[1800]);
assign l_36[740]    = ( l_37 [950] & !i[1800]) | ( l_37 [951] &  i[1800]);
assign l_36[741]    = ( l_37 [952] & !i[1800]) | ( l_37 [953] &  i[1800]);
assign l_36[742]    = ( l_37 [954] & !i[1800]) | ( l_37 [955] &  i[1800]);
assign l_36[743]    = ( l_37 [956] & !i[1800]) | ( l_37 [957] &  i[1800]);
assign l_36[744]    = ( l_37 [958] & !i[1800]) | ( l_37 [959] &  i[1800]);
assign l_36[745]    = ( l_37 [960] & !i[1800]) | ( l_37 [961] &  i[1800]);
assign l_36[746]    = ( l_37 [962] & !i[1800]) | ( l_37 [963] &  i[1800]);
assign l_36[747]    = ( l_37 [964] & !i[1800]) | ( l_37 [965] &  i[1800]);
assign l_36[748]    = ( l_37 [966] & !i[1800]) | ( l_37 [967] &  i[1800]);
assign l_36[749]    = ( l_37 [968] & !i[1800]) | ( l_37 [969] &  i[1800]);
assign l_36[750]    = ( l_37 [970] & !i[1800]) | ( l_37 [971] &  i[1800]);
assign l_36[751]    = ( l_37 [972] & !i[1800]) | ( l_37 [973] &  i[1800]);
assign l_36[752]    = ( l_37 [974] & !i[1800]) | ( l_37 [975] &  i[1800]);
assign l_36[753]    = ( l_37 [976] & !i[1800]) | ( l_37 [977] &  i[1800]);
assign l_36[754]    = ( l_37 [978] & !i[1800]) | ( l_37 [979] &  i[1800]);
assign l_36[755]    = ( l_37 [980] & !i[1800]) | ( l_37 [981] &  i[1800]);
assign l_36[756]    = ( l_37 [982] & !i[1800]) | ( l_37 [983] &  i[1800]);
assign l_36[757]    = ( l_37 [984] & !i[1800]) | ( l_37 [985] &  i[1800]);
assign l_36[758]    = ( l_37 [986] & !i[1800]) | ( l_37 [987] &  i[1800]);
assign l_36[759]    = ( l_37 [988] & !i[1800]) | ( l_37 [989] &  i[1800]);
assign l_36[760]    = ( l_37 [990] & !i[1800]) | ( l_37 [991] &  i[1800]);
assign l_36[761]    = ( l_37 [992] & !i[1800]) | ( l_37 [993] &  i[1800]);
assign l_36[762]    = ( l_37 [994] & !i[1800]) | ( l_37 [995] &  i[1800]);
assign l_36[763]    = ( l_37 [996] & !i[1800]) | ( l_37 [997] &  i[1800]);
assign l_36[764]    = ( l_37 [998] & !i[1800]) | ( l_37 [999] &  i[1800]);
assign l_36[765]    = ( l_37 [1000] & !i[1800]) | ( l_37 [1001] &  i[1800]);
assign l_36[766]    = ( l_37 [1002] & !i[1800]) | ( l_37 [1003] &  i[1800]);
assign l_36[767]    = ( l_37 [1004] & !i[1800]) | ( l_37 [1005] &  i[1800]);
assign l_36[768]    = ( l_37 [1006] & !i[1800]) | ( l_37 [1007] &  i[1800]);
assign l_36[769]    = ( l_37 [1008] & !i[1800]) | ( l_37 [1009] &  i[1800]);
assign l_36[770]    = ( l_37 [1010] & !i[1800]) | ( l_37 [1011] &  i[1800]);
assign l_36[771]    = ( l_37 [1012] & !i[1800]) | ( l_37 [1013] &  i[1800]);
assign l_36[772]    = ( l_37 [1014] & !i[1800]) | ( l_37 [1015] &  i[1800]);
assign l_36[773]    = ( l_37 [1016] & !i[1800]) | ( l_37 [1017] &  i[1800]);
assign l_36[774]    = ( l_37 [1018] & !i[1800]) | ( l_37 [1019] &  i[1800]);
assign l_36[775]    = ( l_37 [1020] & !i[1800]) | ( l_37 [1021] &  i[1800]);
assign l_36[776]    = ( l_37 [1022] & !i[1800]) | ( l_37 [1023] &  i[1800]);
assign l_36[777]    = ( l_37 [1024] & !i[1800]) | ( l_37 [1025] &  i[1800]);
assign l_36[778]    = ( l_37 [1026] & !i[1800]) | ( l_37 [1027] &  i[1800]);
assign l_36[779]    = ( l_37 [1028] & !i[1800]) | ( l_37 [1029] &  i[1800]);
assign l_36[780]    = ( l_37 [1030] & !i[1800]) | ( l_37 [1031] &  i[1800]);
assign l_36[781]    = ( l_37 [1032] & !i[1800]) | ( l_37 [1033] &  i[1800]);
assign l_36[782]    = ( l_37 [1034] & !i[1800]) | ( l_37 [1035] &  i[1800]);
assign l_36[783]    = ( l_37 [1036] & !i[1800]) | ( l_37 [1037] &  i[1800]);
assign l_36[784]    = ( l_37 [1038] & !i[1800]) | ( l_37 [1039] &  i[1800]);
assign l_36[785]    = ( l_37 [1040] & !i[1800]) | ( l_37 [1041] &  i[1800]);
assign l_36[786]    = ( l_37 [1042] & !i[1800]) | ( l_37 [1043] &  i[1800]);
assign l_36[787]    = ( l_37 [1044] & !i[1800]) | ( l_37 [1045] &  i[1800]);
assign l_36[788]    = ( l_37 [1046] & !i[1800]) | ( l_37 [1047] &  i[1800]);
assign l_36[789]    = ( l_37 [1048] & !i[1800]) | ( l_37 [1049] &  i[1800]);
assign l_36[790]    = ( l_37 [1050] & !i[1800]) | ( l_37 [1051] &  i[1800]);
assign l_36[791]    = ( l_37 [1052] & !i[1800]) | ( l_37 [1053] &  i[1800]);
assign l_36[792]    = ( l_37 [1054] & !i[1800]) | ( l_37 [1055] &  i[1800]);
assign l_36[793]    = ( l_37 [1056] & !i[1800]) | ( l_37 [1057] &  i[1800]);
assign l_36[794]    = ( l_37 [1058] & !i[1800]) | ( l_37 [1059] &  i[1800]);
assign l_36[795]    = ( l_37 [1060] & !i[1800]) | ( l_37 [1061] &  i[1800]);
assign l_36[796]    = ( l_37 [1062] & !i[1800]) | ( l_37 [1063] &  i[1800]);
assign l_36[797]    = ( l_37 [1064] & !i[1800]) | ( l_37 [1065] &  i[1800]);
assign l_36[798]    = ( l_37 [1066] & !i[1800]) | ( l_37 [1067] &  i[1800]);
assign l_36[799]    = ( l_37 [1068] & !i[1800]) | ( l_37 [1069] &  i[1800]);
assign l_36[800]    = ( l_37 [1070] & !i[1800]) | ( l_37 [1071] &  i[1800]);
assign l_36[801]    = ( l_37 [1072] & !i[1800]) | ( l_37 [1073] &  i[1800]);
assign l_36[802]    = ( l_37 [1074] & !i[1800]) | ( l_37 [1075] &  i[1800]);
assign l_36[803]    = ( l_37 [1076] & !i[1800]) | ( l_37 [1077] &  i[1800]);
assign l_36[804]    = ( l_37 [1078] & !i[1800]) | ( l_37 [1079] &  i[1800]);
assign l_36[805]    = ( l_37 [1080] & !i[1800]) | ( l_37 [1081] &  i[1800]);
assign l_36[806]    = ( l_37 [1082] & !i[1800]) | ( l_37 [1083] &  i[1800]);
assign l_36[807]    = ( l_37 [1084] & !i[1800]) | ( l_37 [1085] &  i[1800]);
assign l_36[808]    = ( l_37 [1086] & !i[1800]) | ( l_37 [1087] &  i[1800]);
assign l_36[809]    = ( l_37 [1088] & !i[1800]) | ( l_37 [1089] &  i[1800]);
assign l_36[810]    = ( l_37 [1090] & !i[1800]) | ( l_37 [1091] &  i[1800]);
assign l_36[811]    = ( l_37 [1092] & !i[1800]) | ( l_37 [1093] &  i[1800]);
assign l_36[812]    = ( l_37 [1094] & !i[1800]) | ( l_37 [1095] &  i[1800]);
assign l_36[813]    = ( l_37 [1096] & !i[1800]) | ( l_37 [1097] &  i[1800]);
assign l_36[814]    = ( l_37 [1098] & !i[1800]) | ( l_37 [1099] &  i[1800]);
assign l_36[815]    = ( l_37 [1100] & !i[1800]) | ( l_37 [1101] &  i[1800]);
assign l_36[816]    = ( l_37 [1102] & !i[1800]) | ( l_37 [1103] &  i[1800]);
assign l_36[817]    = ( l_37 [1104] & !i[1800]) | ( l_37 [1105] &  i[1800]);
assign l_36[818]    = ( l_37 [1106] & !i[1800]) | ( l_37 [1107] &  i[1800]);
assign l_36[819]    = ( l_37 [1108] & !i[1800]) | ( l_37 [1109] &  i[1800]);
assign l_36[820]    = ( l_37 [1110] & !i[1800]) | ( l_37 [1111] &  i[1800]);
assign l_36[821]    = ( l_37 [1112] & !i[1800]) | ( l_37 [1113] &  i[1800]);
assign l_36[822]    = ( l_37 [1114] & !i[1800]) | ( l_37 [1115] &  i[1800]);
assign l_36[823]    = ( l_37 [1116] & !i[1800]) | ( l_37 [1117] &  i[1800]);
assign l_36[824]    = ( l_37 [1118] & !i[1800]) | ( l_37 [1119] &  i[1800]);
assign l_36[825]    = ( l_37 [1120] & !i[1800]) | ( l_37 [1121] &  i[1800]);
assign l_36[826]    = ( l_37 [1122] & !i[1800]) | ( l_37 [1123] &  i[1800]);
assign l_36[827]    = ( l_37 [1124] & !i[1800]) | ( l_37 [1125] &  i[1800]);
assign l_36[828]    = ( l_37 [1126] & !i[1800]) | ( l_37 [1127] &  i[1800]);
assign l_36[829]    = ( l_37 [1128] & !i[1800]) | ( l_37 [1129] &  i[1800]);
assign l_36[830]    = ( l_37 [1130] & !i[1800]) | ( l_37 [1131] &  i[1800]);
assign l_36[831]    = ( l_37 [1132] & !i[1800]) | ( l_37 [1133] &  i[1800]);
assign l_36[832]    = ( l_37 [1134] & !i[1800]) | ( l_37 [1135] &  i[1800]);
assign l_36[833]    = ( l_37 [1136] & !i[1800]) | ( l_37 [1137] &  i[1800]);
assign l_36[834]    = ( l_37 [1138] & !i[1800]) | ( l_37 [1139] &  i[1800]);
assign l_36[835]    = ( l_37 [1140] & !i[1800]) | ( l_37 [1141] &  i[1800]);
assign l_36[836]    = ( l_37 [1142] & !i[1800]) | ( l_37 [1143] &  i[1800]);
assign l_36[837]    = ( l_37 [1144] & !i[1800]) | ( l_37 [1145] &  i[1800]);
assign l_36[838]    = ( l_37 [1146] & !i[1800]) | ( l_37 [1147] &  i[1800]);
assign l_36[839]    = ( l_37 [1148] & !i[1800]) | ( l_37 [1149] &  i[1800]);
assign l_36[840]    = ( l_37 [1150] & !i[1800]) | ( l_37 [1151] &  i[1800]);
assign l_36[841]    = ( l_37 [1152] & !i[1800]) | ( l_37 [1153] &  i[1800]);
assign l_36[842]    = ( l_37 [1154] & !i[1800]) | ( l_37 [1155] &  i[1800]);
assign l_36[843]    = ( l_37 [1156] & !i[1800]) | ( l_37 [1157] &  i[1800]);
assign l_36[844]    = ( l_37 [1158] & !i[1800]) | ( l_37 [1159] &  i[1800]);
assign l_36[845]    = ( l_37 [1160] & !i[1800]) | ( l_37 [1161] &  i[1800]);
assign l_36[846]    = ( l_37 [1162] & !i[1800]) | ( l_37 [1163] &  i[1800]);
assign l_36[847]    = ( l_37 [1164] & !i[1800]) | ( l_37 [1165] &  i[1800]);
assign l_36[848]    = ( l_37 [1166] & !i[1800]) | ( l_37 [1167] &  i[1800]);
assign l_36[849]    = ( l_37 [1168] & !i[1800]) | ( l_37 [1169] &  i[1800]);
assign l_36[850]    = ( l_37 [1170] & !i[1800]) | ( l_37 [1171] &  i[1800]);
assign l_36[851]    = ( l_37 [1172] & !i[1800]) | ( l_37 [1173] &  i[1800]);
assign l_36[852]    = ( l_37 [1174] & !i[1800]) | ( l_37 [1175] &  i[1800]);
assign l_36[853]    = ( l_37 [1176] & !i[1800]) | ( l_37 [1177] &  i[1800]);
assign l_36[854]    = ( l_37 [1178] & !i[1800]) | ( l_37 [1179] &  i[1800]);
assign l_36[855]    = ( l_37 [1180] & !i[1800]) | ( l_37 [1181] &  i[1800]);
assign l_36[856]    = ( l_37 [1182] & !i[1800]) | ( l_37 [1183] &  i[1800]);
assign l_36[857]    = ( l_37 [1184] & !i[1800]) | ( l_37 [1185] &  i[1800]);
assign l_36[858]    = ( l_37 [1186] & !i[1800]) | ( l_37 [1187] &  i[1800]);
assign l_36[859]    = ( l_37 [1188] & !i[1800]) | ( l_37 [1189] &  i[1800]);
assign l_36[860]    = ( l_37 [1190] & !i[1800]) | ( l_37 [1191] &  i[1800]);
assign l_36[861]    = ( l_37 [1192] & !i[1800]) | ( l_37 [1193] &  i[1800]);
assign l_36[862]    = ( l_37 [1194] & !i[1800]) | ( l_37 [1195] &  i[1800]);
assign l_36[863]    = ( l_37 [1196] & !i[1800]) | ( l_37 [1197] &  i[1800]);
assign l_36[864]    = ( l_37 [1198] & !i[1800]) | ( l_37 [1199] &  i[1800]);
assign l_36[865]    = ( l_37 [1200] & !i[1800]) | ( l_37 [1201] &  i[1800]);
assign l_36[866]    = ( l_37 [1202] & !i[1800]) | ( l_37 [1203] &  i[1800]);
assign l_36[867]    = ( l_37 [1204] & !i[1800]) | ( l_37 [1205] &  i[1800]);
assign l_36[868]    = ( l_37 [1206] & !i[1800]) | ( l_37 [1207] &  i[1800]);
assign l_36[869]    = ( l_37 [1208] & !i[1800]) | ( l_37 [1209] &  i[1800]);
assign l_36[870]    = ( l_37 [1210] & !i[1800]) | ( l_37 [1211] &  i[1800]);
assign l_36[871]    = ( l_37 [1212] & !i[1800]) | ( l_37 [1213] &  i[1800]);
assign l_36[872]    = ( l_37 [1214] & !i[1800]) | ( l_37 [1215] &  i[1800]);
assign l_36[873]    = ( l_37 [1216] & !i[1800]) | ( l_37 [1217] &  i[1800]);
assign l_36[874]    = ( l_37 [1218] & !i[1800]) | ( l_37 [1219] &  i[1800]);
assign l_36[875]    = ( l_37 [1220] & !i[1800]) | ( l_37 [1221] &  i[1800]);
assign l_36[876]    = ( l_37 [1222] & !i[1800]) | ( l_37 [1223] &  i[1800]);
assign l_36[877]    = ( l_37 [1224] & !i[1800]) | ( l_37 [1225] &  i[1800]);
assign l_36[878]    = ( l_37 [1226] & !i[1800]) | ( l_37 [1227] &  i[1800]);
assign l_36[879]    = ( l_37 [1228] & !i[1800]) | ( l_37 [1229] &  i[1800]);
assign l_36[880]    = ( l_37 [1230] & !i[1800]) | ( l_37 [1231] &  i[1800]);
assign l_36[881]    = ( l_37 [1232] & !i[1800]) | ( l_37 [1233] &  i[1800]);
assign l_36[882]    = ( l_37 [1234] & !i[1800]) | ( l_37 [1235] &  i[1800]);
assign l_36[883]    = ( l_37 [1236] & !i[1800]) | ( l_37 [1237] &  i[1800]);
assign l_36[884]    = ( l_37 [1238] & !i[1800]) | ( l_37 [1239] &  i[1800]);
assign l_36[885]    = ( l_37 [1240] & !i[1800]) | ( l_37 [1241] &  i[1800]);
assign l_36[886]    = ( l_37 [1242] & !i[1800]) | ( l_37 [1243] &  i[1800]);
assign l_36[887]    = ( l_37 [1244] & !i[1800]) | ( l_37 [1245] &  i[1800]);
assign l_36[888]    = ( l_37 [1246] & !i[1800]) | ( l_37 [1247] &  i[1800]);
assign l_36[889]    = ( l_37 [1248] & !i[1800]) | ( l_37 [1249] &  i[1800]);
assign l_36[890]    = ( l_37 [1250] & !i[1800]) | ( l_37 [1251] &  i[1800]);
assign l_36[891]    = ( l_37 [1252] & !i[1800]) | ( l_37 [1253] &  i[1800]);
assign l_36[892]    = ( l_37 [1254] & !i[1800]) | ( l_37 [1255] &  i[1800]);
assign l_36[893]    = ( l_37 [1256] & !i[1800]) | ( l_37 [1257] &  i[1800]);
assign l_36[894]    = ( l_37 [1258] & !i[1800]) | ( l_37 [1259] &  i[1800]);
assign l_36[895]    = ( l_37 [1260] & !i[1800]) | ( l_37 [1261] &  i[1800]);
assign l_36[896]    = ( l_37 [1262] & !i[1800]) | ( l_37 [1263] &  i[1800]);
assign l_36[897]    = ( l_37 [1264] & !i[1800]) | ( l_37 [1265] &  i[1800]);
assign l_36[898]    = ( l_37 [1266] & !i[1800]) | ( l_37 [1267] &  i[1800]);
assign l_36[899]    = ( l_37 [1268] & !i[1800]) | ( l_37 [1269] &  i[1800]);
assign l_36[900]    = ( l_37 [1270] & !i[1800]) | ( l_37 [1271] &  i[1800]);
assign l_36[901]    = ( l_37 [1272] & !i[1800]) | ( l_37 [1273] &  i[1800]);
assign l_36[902]    = ( l_37 [1274] & !i[1800]) | ( l_37 [1275] &  i[1800]);
assign l_36[903]    = ( l_37 [1276] & !i[1800]) | ( l_37 [1277] &  i[1800]);
assign l_36[904]    = ( l_37 [1278] & !i[1800]) | ( l_37 [1279] &  i[1800]);
assign l_36[905]    = ( l_37 [1280] & !i[1800]) | ( l_37 [1281] &  i[1800]);
assign l_36[906]    = ( l_37 [1282] & !i[1800]) | ( l_37 [1283] &  i[1800]);
assign l_36[907]    = ( l_37 [1284] & !i[1800]) | ( l_37 [1285] &  i[1800]);
assign l_36[908]    = ( l_37 [1286] & !i[1800]) | ( l_37 [1287] &  i[1800]);
assign l_36[909]    = ( l_37 [1288] & !i[1800]) | ( l_37 [1289] &  i[1800]);
assign l_36[910]    = ( l_37 [1290] & !i[1800]) | ( l_37 [1291] &  i[1800]);
assign l_36[911]    = ( l_37 [1292] & !i[1800]) | ( l_37 [1293] &  i[1800]);
assign l_36[912]    = ( l_37 [1294] & !i[1800]) | ( l_37 [1295] &  i[1800]);
assign l_36[913]    = ( l_37 [1296] & !i[1800]) | ( l_37 [1297] &  i[1800]);
assign l_36[914]    = ( l_37 [1298] & !i[1800]) | ( l_37 [1299] &  i[1800]);
assign l_36[915]    = ( l_37 [1300] & !i[1800]) | ( l_37 [1301] &  i[1800]);
assign l_36[916]    = ( l_37 [1302] & !i[1800]) | ( l_37 [1303] &  i[1800]);
assign l_36[917]    = ( l_37 [1304] & !i[1800]) | ( l_37 [1305] &  i[1800]);
assign l_36[918]    = ( l_37 [1306] & !i[1800]) | ( l_37 [1307] &  i[1800]);
assign l_36[919]    = ( l_37 [1308] & !i[1800]) | ( l_37 [1309] &  i[1800]);
assign l_36[920]    = ( l_37 [1310] & !i[1800]) | ( l_37 [1311] &  i[1800]);
assign l_36[921]    = ( l_37 [1312] & !i[1800]) | ( l_37 [1313] &  i[1800]);
assign l_36[922]    = ( l_37 [1314] & !i[1800]) | ( l_37 [1315] &  i[1800]);
assign l_36[923]    = ( l_37 [1316] & !i[1800]) | ( l_37 [1317] &  i[1800]);
assign l_36[924]    = ( l_37 [1318] & !i[1800]) | ( l_37 [1319] &  i[1800]);
assign l_36[925]    = ( l_37 [1320] & !i[1800]) | ( l_37 [1321] &  i[1800]);
assign l_36[926]    = ( l_37 [1322] & !i[1800]) | ( l_37 [1323] &  i[1800]);
assign l_36[927]    = ( l_37 [1324] & !i[1800]) | ( l_37 [1325] &  i[1800]);
assign l_36[928]    = ( l_37 [1326] & !i[1800]) | ( l_37 [1327] &  i[1800]);
assign l_36[929]    = ( l_37 [1328] & !i[1800]) | ( l_37 [1329] &  i[1800]);
assign l_36[930]    = ( l_37 [1330] & !i[1800]) | ( l_37 [1331] &  i[1800]);
assign l_36[931]    = ( l_37 [1332] & !i[1800]) | ( l_37 [1333] &  i[1800]);
assign l_36[932]    = ( l_37 [1334] & !i[1800]) | ( l_37 [1335] &  i[1800]);
assign l_36[933]    = ( l_37 [1336] & !i[1800]) | ( l_37 [1337] &  i[1800]);
assign l_36[934]    = ( l_37 [1338] & !i[1800]) | ( l_37 [1339] &  i[1800]);
assign l_36[935]    = ( l_37 [1340] & !i[1800]) | ( l_37 [1341] &  i[1800]);
assign l_36[936]    = ( l_37 [1342] & !i[1800]) | ( l_37 [1343] &  i[1800]);
assign l_36[937]    = ( l_37 [1344] & !i[1800]) | ( l_37 [1345] &  i[1800]);
assign l_36[938]    = ( l_37 [1346] & !i[1800]) | ( l_37 [1347] &  i[1800]);
assign l_36[939]    = ( l_37 [1348] & !i[1800]) | ( l_37 [1349] &  i[1800]);
assign l_36[940]    = ( l_37 [1350] & !i[1800]) | ( l_37 [1351] &  i[1800]);
assign l_36[941]    = ( l_37 [1352] & !i[1800]) | ( l_37 [1353] &  i[1800]);
assign l_36[942]    = ( l_37 [1354] & !i[1800]) | ( l_37 [1355] &  i[1800]);
assign l_36[943]    = ( l_37 [1356] & !i[1800]) | ( l_37 [1357] &  i[1800]);
assign l_36[944]    = ( l_37 [1358] & !i[1800]) | ( l_37 [1359] &  i[1800]);
assign l_36[945]    = ( l_37 [1360] & !i[1800]) | ( l_37 [1361] &  i[1800]);
assign l_36[946]    = ( l_37 [1362] & !i[1800]) | ( l_37 [1363] &  i[1800]);
assign l_36[947]    = ( l_37 [1364] & !i[1800]) | ( l_37 [1365] &  i[1800]);
assign l_36[948]    = ( l_37 [1366] & !i[1800]) | ( l_37 [1367] &  i[1800]);
assign l_36[949]    = ( l_37 [1368] & !i[1800]) | ( l_37 [1369] &  i[1800]);
assign l_36[950]    = ( l_37 [1370] & !i[1800]) | ( l_37 [1371] &  i[1800]);
assign l_36[951]    = ( l_37 [1372] & !i[1800]) | ( l_37 [1373] &  i[1800]);
assign l_36[952]    = ( l_37 [1374] & !i[1800]) | ( l_37 [1375] &  i[1800]);
assign l_36[953]    = ( l_37 [1376] & !i[1800]) | ( l_37 [1377] &  i[1800]);
assign l_36[954]    = ( l_37 [1378] & !i[1800]) | ( l_37 [1379] &  i[1800]);
assign l_36[955]    = ( l_37 [1380] & !i[1800]) | ( l_37 [1381] &  i[1800]);
assign l_36[956]    = ( l_37 [1382] & !i[1800]) | ( l_37 [1383] &  i[1800]);
assign l_36[957]    = ( l_37 [1384] & !i[1800]) | ( l_37 [1385] &  i[1800]);
assign l_36[958]    = ( l_37 [1386] & !i[1800]) | ( l_37 [1387] &  i[1800]);
assign l_36[959]    = ( l_37 [1388] & !i[1800]) | ( l_37 [1389] &  i[1800]);
assign l_36[960]    = ( l_37 [1390] & !i[1800]) | ( l_37 [1391] &  i[1800]);
assign l_36[961]    = ( l_37 [1392] & !i[1800]) | ( l_37 [1393] &  i[1800]);
assign l_36[962]    = ( l_37 [1394] & !i[1800]) | ( l_37 [1395] &  i[1800]);
assign l_36[963]    = ( l_37 [1396] & !i[1800]) | ( l_37 [1397] &  i[1800]);
assign l_36[964]    = ( l_37 [1398] & !i[1800]) | ( l_37 [1399] &  i[1800]);
assign l_36[965]    = ( l_37 [1400] & !i[1800]) | ( l_37 [1401] &  i[1800]);
assign l_36[966]    = ( l_37 [1402] & !i[1800]) | ( l_37 [1403] &  i[1800]);
assign l_36[967]    = ( l_37 [1404] & !i[1800]) | ( l_37 [1405] &  i[1800]);
assign l_36[968]    = ( l_37 [1406] & !i[1800]) | ( l_37 [1407] &  i[1800]);
assign l_36[969]    = ( l_37 [1408] & !i[1800]) | ( l_37 [1409] &  i[1800]);
assign l_36[970]    = ( l_37 [1410] & !i[1800]) | ( l_37 [1411] &  i[1800]);
assign l_36[971]    = ( l_37 [1412] & !i[1800]) | ( l_37 [1413] &  i[1800]);
assign l_36[972]    = ( l_37 [1414] & !i[1800]) | ( l_37 [1415] &  i[1800]);
assign l_36[973]    = ( l_37 [1416] & !i[1800]) | ( l_37 [1417] &  i[1800]);
assign l_36[974]    = ( l_37 [1418] & !i[1800]) | ( l_37 [1419] &  i[1800]);
assign l_36[975]    = ( l_37 [1420] & !i[1800]) | ( l_37 [1421] &  i[1800]);
assign l_36[976]    = ( l_37 [1422] & !i[1800]) | ( l_37 [1423] &  i[1800]);
assign l_36[977]    = ( l_37 [1424] & !i[1800]) | ( l_37 [1425] &  i[1800]);
assign l_36[978]    = ( l_37 [1426] & !i[1800]) | ( l_37 [1427] &  i[1800]);
assign l_36[979]    = ( l_37 [1428] & !i[1800]) | ( l_37 [1429] &  i[1800]);
assign l_36[980]    = ( l_37 [1430] & !i[1800]) | ( l_37 [1431] &  i[1800]);
assign l_36[981]    = ( l_37 [1432] & !i[1800]) | ( l_37 [1433] &  i[1800]);
assign l_36[982]    = ( l_37 [1434] & !i[1800]) | ( l_37 [1435] &  i[1800]);
assign l_36[983]    = ( l_37 [1436] & !i[1800]) | ( l_37 [1437] &  i[1800]);
assign l_36[984]    = ( l_37 [1438] & !i[1800]) | ( l_37 [1439] &  i[1800]);
assign l_36[985]    = ( l_37 [1440] & !i[1800]) | ( l_37 [1441] &  i[1800]);
assign l_36[986]    = ( l_37 [1442] & !i[1800]) | ( l_37 [1443] &  i[1800]);
assign l_36[987]    = ( l_37 [1444] & !i[1800]) | ( l_37 [1445] &  i[1800]);
assign l_36[988]    = ( l_37 [1446] & !i[1800]) | ( l_37 [1447] &  i[1800]);
assign l_36[989]    = ( l_37 [1448] & !i[1800]) | ( l_37 [1449] &  i[1800]);
assign l_36[990]    = ( l_37 [1450] & !i[1800]) | ( l_37 [1451] &  i[1800]);
assign l_36[991]    = ( l_37 [1452] & !i[1800]) | ( l_37 [1453] &  i[1800]);
assign l_36[992]    = ( l_37 [1454] & !i[1800]) | ( l_37 [1455] &  i[1800]);
assign l_36[993]    = ( l_37 [1456] & !i[1800]) | ( l_37 [1457] &  i[1800]);
assign l_36[994]    = ( l_37 [1458] & !i[1800]) | ( l_37 [1459] &  i[1800]);
assign l_36[995]    = ( l_37 [1460] & !i[1800]) | ( l_37 [1461] &  i[1800]);
assign l_36[996]    = ( l_37 [1462] & !i[1800]) | ( l_37 [1463] &  i[1800]);
assign l_36[997]    = ( l_37 [1464] & !i[1800]) | ( l_37 [1465] &  i[1800]);
assign l_36[998]    = ( l_37 [1466] & !i[1800]) | ( l_37 [1467] &  i[1800]);
assign l_36[999]    = ( l_37 [1468] & !i[1800]) | ( l_37 [1469] &  i[1800]);
assign l_36[1000]    = ( l_37 [1470] & !i[1800]) | ( l_37 [1471] &  i[1800]);
assign l_36[1001]    = ( l_37 [1472] & !i[1800]) | ( l_37 [1473] &  i[1800]);
assign l_36[1002]    = ( l_37 [1474] & !i[1800]) | ( l_37 [1475] &  i[1800]);
assign l_36[1003]    = ( l_37 [1476] & !i[1800]) | ( l_37 [1477] &  i[1800]);
assign l_36[1004]    = ( l_37 [1478] & !i[1800]) | ( l_37 [1479] &  i[1800]);
assign l_36[1005]    = ( l_37 [1480] & !i[1800]) | ( l_37 [1481] &  i[1800]);
assign l_36[1006]    = ( l_37 [1482] & !i[1800]) | ( l_37 [1483] &  i[1800]);
assign l_36[1007]    = ( l_37 [1484] & !i[1800]) | ( l_37 [1485] &  i[1800]);
assign l_36[1008]    = ( l_37 [1486] & !i[1800]) | ( l_37 [1487] &  i[1800]);
assign l_36[1009]    = ( l_37 [1488] & !i[1800]) | ( l_37 [1489] &  i[1800]);
assign l_36[1010]    = ( l_37 [1490] & !i[1800]) | ( l_37 [1491] &  i[1800]);
assign l_36[1011]    = ( l_37 [1492] & !i[1800]) | ( l_37 [1493] &  i[1800]);
assign l_36[1012]    = ( l_37 [1494] & !i[1800]) | ( l_37 [1495] &  i[1800]);
assign l_36[1013]    = ( l_37 [1496] & !i[1800]) | ( l_37 [1497] &  i[1800]);
assign l_36[1014]    = ( l_37 [1498] & !i[1800]) | ( l_37 [1499] &  i[1800]);
assign l_36[1015]    = ( l_37 [1500] & !i[1800]) | ( l_37 [1501] &  i[1800]);
assign l_36[1016]    = ( l_37 [1502] & !i[1800]) | ( l_37 [1503] &  i[1800]);
assign l_36[1017]    = ( l_37 [1504] & !i[1800]) | ( l_37 [1505] &  i[1800]);
assign l_36[1018]    = ( l_37 [1506] & !i[1800]) | ( l_37 [1507] &  i[1800]);
assign l_36[1019]    = ( l_37 [1508] & !i[1800]) | ( l_37 [1509] &  i[1800]);
assign l_36[1020]    = ( l_37 [1510] & !i[1800]) | ( l_37 [1511] &  i[1800]);
assign l_36[1021]    = ( l_37 [1512] & !i[1800]) | ( l_37 [1513] &  i[1800]);
assign l_36[1022]    = ( l_37 [1514] & !i[1800]) | ( l_37 [1515] &  i[1800]);
assign l_36[1023]    = ( l_37 [1516] & !i[1800]) | ( l_37 [1517] &  i[1800]);
assign l_36[1024]    = ( l_37 [1518] & !i[1800]) | ( l_37 [1519] &  i[1800]);
assign l_36[1025]    = ( l_37 [1520] & !i[1800]) | ( l_37 [1521] &  i[1800]);
assign l_36[1026]    = ( l_37 [1522] & !i[1800]) | ( l_37 [1523] &  i[1800]);
assign l_36[1027]    = ( l_37 [1524] & !i[1800]) | ( l_37 [1525] &  i[1800]);
assign l_36[1028]    = ( l_37 [1526] & !i[1800]) | ( l_37 [1527] &  i[1800]);
assign l_36[1029]    = ( l_37 [1528] & !i[1800]) | ( l_37 [1529] &  i[1800]);
assign l_36[1030]    = ( l_37 [1530] & !i[1800]) | ( l_37 [1531] &  i[1800]);
assign l_36[1031]    = ( l_37 [1532] & !i[1800]) | ( l_37 [1533] &  i[1800]);
assign l_36[1032]    = ( l_37 [1534] & !i[1800]) | ( l_37 [1535] &  i[1800]);
assign l_36[1033]    = ( l_37 [1536] & !i[1800]) | ( l_37 [1537] &  i[1800]);
assign l_36[1034]    = ( l_37 [1538] & !i[1800]) | ( l_37 [1539] &  i[1800]);
assign l_36[1035]    = ( l_37 [1540] & !i[1800]) | ( l_37 [1541] &  i[1800]);
assign l_36[1036]    = ( l_37 [1542] & !i[1800]) | ( l_37 [1543] &  i[1800]);
assign l_36[1037]    = ( l_37 [1544] & !i[1800]) | ( l_37 [1545] &  i[1800]);
assign l_36[1038]    = ( l_37 [1546] & !i[1800]) | ( l_37 [1547] &  i[1800]);
assign l_36[1039]    = ( l_37 [1548] & !i[1800]) | ( l_37 [1549] &  i[1800]);
assign l_36[1040]    = ( l_37 [1550] & !i[1800]) | ( l_37 [1551] &  i[1800]);
assign l_36[1041]    = ( l_37 [1552] & !i[1800]) | ( l_37 [1553] &  i[1800]);
assign l_37[0]    = ( l_38 [0]);
assign l_37[1]    = ( l_38 [1] & !i[1815]);
assign l_37[2]    = ( l_38 [2] & !i[1815]);
assign l_37[3]    = (!i[1815]) | ( l_38 [3] &  i[1815]);
assign l_37[4]    = (!i[1815]) | ( l_38 [4] &  i[1815]);
assign l_37[5]    = ( l_38 [5] & !i[1815]);
assign l_37[6]    = ( l_38 [6] & !i[1815]);
assign l_37[7]    = (!i[1815]) | ( l_38 [7] &  i[1815]);
assign l_37[8]    = (!i[1815]) | ( l_38 [8] &  i[1815]);
assign l_37[9]    = ( l_38 [9] & !i[1815]) | ( l_38 [10] &  i[1815]);
assign l_37[10]    = ( l_38 [10]);
assign l_37[11]    = ( l_38 [11] & !i[1815]) | ( l_38 [10] &  i[1815]);
assign l_37[12]    = ( l_38 [10] & !i[1815]) | ( l_38 [12] &  i[1815]);
assign l_37[13]    = ( l_38 [10] & !i[1815]) | ( l_38 [13] &  i[1815]);
assign l_37[14]    = ( l_38 [14] & !i[1815]) | ( l_38 [10] &  i[1815]);
assign l_37[15]    = ( l_38 [15] & !i[1815]) | ( l_38 [10] &  i[1815]);
assign l_37[16]    = ( l_38 [10] & !i[1815]) | ( l_38 [16] &  i[1815]);
assign l_37[17]    = ( l_38 [10] & !i[1815]) | ( l_38 [17] &  i[1815]);
assign l_37[18]    = ( l_38 [18] & !i[1815]) | ( l_38 [19] &  i[1815]);
assign l_37[19]    = ( l_38 [20] & !i[1815]) | ( l_38 [21] &  i[1815]);
assign l_37[20]    = ( l_38 [22] & !i[1815]) | ( l_38 [23] &  i[1815]);
assign l_37[21]    = ( l_38 [24] & !i[1815]) | ( l_38 [25] &  i[1815]);
assign l_37[22]    = ( l_38 [26] & !i[1815]) | ( l_38 [27] &  i[1815]);
assign l_37[23]    = ( l_38 [28] & !i[1815]) | ( l_38 [29] &  i[1815]);
assign l_37[24]    = ( l_38 [30] & !i[1815]) | ( l_38 [31] &  i[1815]);
assign l_37[25]    = ( l_38 [32] & !i[1815]) | ( l_38 [33] &  i[1815]);
assign l_37[26]    = ( l_38 [34] & !i[1815]) | ( l_38 [35] &  i[1815]);
assign l_37[27]    = ( l_38 [36] & !i[1815]) | ( l_38 [37] &  i[1815]);
assign l_37[28]    = ( l_38 [38] & !i[1815]) | ( l_38 [39] &  i[1815]);
assign l_37[29]    = ( l_38 [40] & !i[1815]) | ( l_38 [41] &  i[1815]);
assign l_37[30]    = ( l_38 [42] & !i[1815]) | ( l_38 [43] &  i[1815]);
assign l_37[31]    = ( l_38 [44] & !i[1815]) | ( l_38 [45] &  i[1815]);
assign l_37[32]    = ( l_38 [46] & !i[1815]) | ( l_38 [47] &  i[1815]);
assign l_37[33]    = ( l_38 [48] & !i[1815]) | ( l_38 [49] &  i[1815]);
assign l_37[34]    = ( l_38 [50] & !i[1815]) | ( l_38 [51] &  i[1815]);
assign l_37[35]    = ( l_38 [52] & !i[1815]) | ( l_38 [53] &  i[1815]);
assign l_37[36]    = ( l_38 [54] & !i[1815]) | ( l_38 [55] &  i[1815]);
assign l_37[37]    = ( l_38 [56] & !i[1815]) | ( l_38 [57] &  i[1815]);
assign l_37[38]    = ( l_38 [58] & !i[1815]) | ( l_38 [59] &  i[1815]);
assign l_37[39]    = ( l_38 [60] & !i[1815]) | ( l_38 [61] &  i[1815]);
assign l_37[40]    = ( l_38 [62] & !i[1815]) | ( l_38 [63] &  i[1815]);
assign l_37[41]    = ( l_38 [64] & !i[1815]) | ( l_38 [65] &  i[1815]);
assign l_37[42]    = ( l_38 [66] & !i[1815]) | ( l_38 [67] &  i[1815]);
assign l_37[43]    = ( l_38 [68] & !i[1815]) | ( l_38 [69] &  i[1815]);
assign l_37[44]    = ( l_38 [70] & !i[1815]) | ( l_38 [71] &  i[1815]);
assign l_37[45]    = ( l_38 [72] & !i[1815]) | ( l_38 [73] &  i[1815]);
assign l_37[46]    = ( l_38 [74] & !i[1815]) | ( l_38 [75] &  i[1815]);
assign l_37[47]    = ( l_38 [76] & !i[1815]) | ( l_38 [77] &  i[1815]);
assign l_37[48]    = ( l_38 [78] & !i[1815]) | ( l_38 [79] &  i[1815]);
assign l_37[49]    = ( l_38 [80] & !i[1815]) | ( l_38 [81] &  i[1815]);
assign l_37[50]    = ( l_38 [82] & !i[1815]) | ( l_38 [83] &  i[1815]);
assign l_37[51]    = ( l_38 [84] & !i[1815]) | ( l_38 [85] &  i[1815]);
assign l_37[52]    = ( l_38 [86] & !i[1815]) | ( l_38 [87] &  i[1815]);
assign l_37[53]    = ( l_38 [88] & !i[1815]) | ( l_38 [89] &  i[1815]);
assign l_37[54]    = ( l_38 [90] & !i[1815]) | ( l_38 [91] &  i[1815]);
assign l_37[55]    = ( l_38 [92] & !i[1815]) | ( l_38 [93] &  i[1815]);
assign l_37[56]    = ( l_38 [94] & !i[1815]) | ( l_38 [95] &  i[1815]);
assign l_37[57]    = ( l_38 [96] & !i[1815]) | ( l_38 [97] &  i[1815]);
assign l_37[58]    = ( l_38 [98] & !i[1815]) | ( l_38 [99] &  i[1815]);
assign l_37[59]    = ( l_38 [100] & !i[1815]) | ( l_38 [101] &  i[1815]);
assign l_37[60]    = ( l_38 [102] & !i[1815]) | ( l_38 [103] &  i[1815]);
assign l_37[61]    = ( l_38 [104] & !i[1815]) | ( l_38 [105] &  i[1815]);
assign l_37[62]    = ( l_38 [106] & !i[1815]) | ( l_38 [107] &  i[1815]);
assign l_37[63]    = ( l_38 [108] & !i[1815]) | ( l_38 [109] &  i[1815]);
assign l_37[64]    = ( l_38 [110] & !i[1815]) | ( l_38 [111] &  i[1815]);
assign l_37[65]    = ( l_38 [112] & !i[1815]) | ( l_38 [113] &  i[1815]);
assign l_37[66]    = ( l_38 [114] & !i[1815]) | ( l_38 [115] &  i[1815]);
assign l_37[67]    = ( l_38 [116] & !i[1815]) | ( l_38 [117] &  i[1815]);
assign l_37[68]    = ( l_38 [118] & !i[1815]) | ( l_38 [119] &  i[1815]);
assign l_37[69]    = ( l_38 [120] & !i[1815]) | ( l_38 [121] &  i[1815]);
assign l_37[70]    = ( l_38 [122] & !i[1815]) | ( l_38 [123] &  i[1815]);
assign l_37[71]    = ( l_38 [124] & !i[1815]) | ( l_38 [125] &  i[1815]);
assign l_37[72]    = ( l_38 [126] & !i[1815]) | ( l_38 [127] &  i[1815]);
assign l_37[73]    = ( l_38 [128] & !i[1815]) | ( l_38 [129] &  i[1815]);
assign l_37[74]    = ( l_38 [130] & !i[1815]) | ( l_38 [131] &  i[1815]);
assign l_37[75]    = ( l_38 [132] & !i[1815]) | ( l_38 [133] &  i[1815]);
assign l_37[76]    = ( l_38 [134] & !i[1815]) | ( l_38 [135] &  i[1815]);
assign l_37[77]    = ( l_38 [136] & !i[1815]) | ( l_38 [137] &  i[1815]);
assign l_37[78]    = ( l_38 [138] & !i[1815]) | ( l_38 [139] &  i[1815]);
assign l_37[79]    = ( l_38 [140] & !i[1815]) | ( l_38 [141] &  i[1815]);
assign l_37[80]    = ( l_38 [142] & !i[1815]) | ( l_38 [143] &  i[1815]);
assign l_37[81]    = ( l_38 [144] & !i[1815]) | ( l_38 [145] &  i[1815]);
assign l_37[82]    = ( l_38 [146] & !i[1815]) | ( l_38 [147] &  i[1815]);
assign l_37[83]    = ( l_38 [148] & !i[1815]) | ( l_38 [149] &  i[1815]);
assign l_37[84]    = ( l_38 [150] & !i[1815]) | ( l_38 [151] &  i[1815]);
assign l_37[85]    = ( l_38 [152] & !i[1815]) | ( l_38 [153] &  i[1815]);
assign l_37[86]    = ( l_38 [154] & !i[1815]) | ( l_38 [155] &  i[1815]);
assign l_37[87]    = ( l_38 [156] & !i[1815]) | ( l_38 [157] &  i[1815]);
assign l_37[88]    = ( l_38 [158] & !i[1815]) | ( l_38 [159] &  i[1815]);
assign l_37[89]    = ( l_38 [160] & !i[1815]) | ( l_38 [161] &  i[1815]);
assign l_37[90]    = ( l_38 [162] & !i[1815]) | ( l_38 [163] &  i[1815]);
assign l_37[91]    = ( l_38 [164] & !i[1815]) | ( l_38 [165] &  i[1815]);
assign l_37[92]    = ( l_38 [166] & !i[1815]) | ( l_38 [167] &  i[1815]);
assign l_37[93]    = ( l_38 [168] & !i[1815]) | ( l_38 [169] &  i[1815]);
assign l_37[94]    = ( l_38 [170] & !i[1815]) | ( l_38 [171] &  i[1815]);
assign l_37[95]    = ( l_38 [172] & !i[1815]) | ( l_38 [173] &  i[1815]);
assign l_37[96]    = ( l_38 [174] & !i[1815]) | ( l_38 [175] &  i[1815]);
assign l_37[97]    = ( l_38 [176] & !i[1815]) | ( l_38 [177] &  i[1815]);
assign l_37[98]    = ( l_38 [178] & !i[1815]) | ( l_38 [179] &  i[1815]);
assign l_37[99]    = ( l_38 [180] & !i[1815]) | ( l_38 [181] &  i[1815]);
assign l_37[100]    = ( l_38 [182] & !i[1815]) | ( l_38 [183] &  i[1815]);
assign l_37[101]    = ( l_38 [184] & !i[1815]) | ( l_38 [185] &  i[1815]);
assign l_37[102]    = ( l_38 [186] & !i[1815]) | ( l_38 [187] &  i[1815]);
assign l_37[103]    = ( l_38 [188] & !i[1815]) | ( l_38 [189] &  i[1815]);
assign l_37[104]    = ( l_38 [190] & !i[1815]) | ( l_38 [191] &  i[1815]);
assign l_37[105]    = ( l_38 [192] & !i[1815]) | ( l_38 [193] &  i[1815]);
assign l_37[106]    = ( l_38 [194] & !i[1815]) | ( l_38 [195] &  i[1815]);
assign l_37[107]    = ( l_38 [196] & !i[1815]) | ( l_38 [197] &  i[1815]);
assign l_37[108]    = ( l_38 [198] & !i[1815]) | ( l_38 [199] &  i[1815]);
assign l_37[109]    = ( l_38 [200] & !i[1815]) | ( l_38 [201] &  i[1815]);
assign l_37[110]    = ( l_38 [202] & !i[1815]) | ( l_38 [203] &  i[1815]);
assign l_37[111]    = ( l_38 [204] & !i[1815]) | ( l_38 [205] &  i[1815]);
assign l_37[112]    = ( l_38 [206] & !i[1815]) | ( l_38 [207] &  i[1815]);
assign l_37[113]    = ( l_38 [208] & !i[1815]) | ( l_38 [209] &  i[1815]);
assign l_37[114]    = ( l_38 [210] & !i[1815]) | ( l_38 [211] &  i[1815]);
assign l_37[115]    = ( l_38 [212] & !i[1815]) | ( l_38 [213] &  i[1815]);
assign l_37[116]    = ( l_38 [214] & !i[1815]) | ( l_38 [215] &  i[1815]);
assign l_37[117]    = ( l_38 [216] & !i[1815]) | ( l_38 [217] &  i[1815]);
assign l_37[118]    = ( l_38 [218] & !i[1815]) | ( l_38 [219] &  i[1815]);
assign l_37[119]    = ( l_38 [220] & !i[1815]) | ( l_38 [221] &  i[1815]);
assign l_37[120]    = ( l_38 [222] & !i[1815]) | ( l_38 [223] &  i[1815]);
assign l_37[121]    = ( l_38 [224] & !i[1815]) | ( l_38 [225] &  i[1815]);
assign l_37[122]    = ( l_38 [226] & !i[1815]) | ( l_38 [227] &  i[1815]);
assign l_37[123]    = ( l_38 [228] & !i[1815]) | ( l_38 [229] &  i[1815]);
assign l_37[124]    = ( l_38 [230] & !i[1815]) | ( l_38 [231] &  i[1815]);
assign l_37[125]    = ( l_38 [232] & !i[1815]) | ( l_38 [233] &  i[1815]);
assign l_37[126]    = ( l_38 [234] & !i[1815]) | ( l_38 [235] &  i[1815]);
assign l_37[127]    = ( l_38 [236] & !i[1815]) | ( l_38 [237] &  i[1815]);
assign l_37[128]    = ( l_38 [238] & !i[1815]) | ( l_38 [239] &  i[1815]);
assign l_37[129]    = ( l_38 [240] & !i[1815]) | ( l_38 [241] &  i[1815]);
assign l_37[130]    = ( l_38 [242] & !i[1815]) | ( l_38 [243] &  i[1815]);
assign l_37[131]    = ( l_38 [244] & !i[1815]) | ( l_38 [245] &  i[1815]);
assign l_37[132]    = ( l_38 [246] & !i[1815]) | ( l_38 [247] &  i[1815]);
assign l_37[133]    = ( l_38 [248] & !i[1815]) | ( l_38 [249] &  i[1815]);
assign l_37[134]    = ( l_38 [250] & !i[1815]) | ( l_38 [251] &  i[1815]);
assign l_37[135]    = ( l_38 [252] & !i[1815]) | ( l_38 [253] &  i[1815]);
assign l_37[136]    = ( l_38 [254] & !i[1815]) | ( l_38 [255] &  i[1815]);
assign l_37[137]    = ( l_38 [256] & !i[1815]) | ( l_38 [257] &  i[1815]);
assign l_37[138]    = ( l_38 [258] & !i[1815]) | ( l_38 [259] &  i[1815]);
assign l_37[139]    = ( l_38 [260] & !i[1815]) | ( l_38 [261] &  i[1815]);
assign l_37[140]    = ( l_38 [262] & !i[1815]) | ( l_38 [263] &  i[1815]);
assign l_37[141]    = ( l_38 [264] & !i[1815]) | ( l_38 [265] &  i[1815]);
assign l_37[142]    = ( l_38 [266] & !i[1815]) | ( l_38 [267] &  i[1815]);
assign l_37[143]    = ( l_38 [268] & !i[1815]) | ( l_38 [269] &  i[1815]);
assign l_37[144]    = ( l_38 [270] & !i[1815]) | ( l_38 [271] &  i[1815]);
assign l_37[145]    = ( l_38 [272] & !i[1815]) | ( l_38 [273] &  i[1815]);
assign l_37[146]    = ( l_38 [274] & !i[1815]) | ( l_38 [275] &  i[1815]);
assign l_37[147]    = ( l_38 [276] & !i[1815]) | ( l_38 [277] &  i[1815]);
assign l_37[148]    = ( l_38 [278] & !i[1815]) | ( l_38 [279] &  i[1815]);
assign l_37[149]    = ( l_38 [280] & !i[1815]) | ( l_38 [281] &  i[1815]);
assign l_37[150]    = ( l_38 [282] & !i[1815]) | ( l_38 [283] &  i[1815]);
assign l_37[151]    = ( l_38 [284] & !i[1815]) | ( l_38 [285] &  i[1815]);
assign l_37[152]    = ( l_38 [286] & !i[1815]) | ( l_38 [287] &  i[1815]);
assign l_37[153]    = ( l_38 [288] & !i[1815]) | ( l_38 [289] &  i[1815]);
assign l_37[154]    = ( l_38 [290] & !i[1815]) | ( l_38 [291] &  i[1815]);
assign l_37[155]    = ( l_38 [292] & !i[1815]) | ( l_38 [293] &  i[1815]);
assign l_37[156]    = ( l_38 [294] & !i[1815]) | ( l_38 [295] &  i[1815]);
assign l_37[157]    = ( l_38 [296] & !i[1815]) | ( l_38 [297] &  i[1815]);
assign l_37[158]    = ( l_38 [298] & !i[1815]) | ( l_38 [299] &  i[1815]);
assign l_37[159]    = ( l_38 [300] & !i[1815]) | ( l_38 [301] &  i[1815]);
assign l_37[160]    = ( l_38 [302] & !i[1815]) | ( l_38 [303] &  i[1815]);
assign l_37[161]    = ( l_38 [304] & !i[1815]) | ( l_38 [305] &  i[1815]);
assign l_37[162]    = ( l_38 [306] & !i[1815]) | ( l_38 [307] &  i[1815]);
assign l_37[163]    = ( l_38 [308] & !i[1815]) | ( l_38 [309] &  i[1815]);
assign l_37[164]    = ( l_38 [310] & !i[1815]) | ( l_38 [311] &  i[1815]);
assign l_37[165]    = ( l_38 [312] & !i[1815]) | ( l_38 [313] &  i[1815]);
assign l_37[166]    = ( l_38 [314] & !i[1815]) | ( l_38 [315] &  i[1815]);
assign l_37[167]    = ( l_38 [316] & !i[1815]) | ( l_38 [317] &  i[1815]);
assign l_37[168]    = ( l_38 [318] & !i[1815]) | ( l_38 [319] &  i[1815]);
assign l_37[169]    = ( l_38 [320] & !i[1815]) | ( l_38 [321] &  i[1815]);
assign l_37[170]    = ( l_38 [322] & !i[1815]) | ( l_38 [323] &  i[1815]);
assign l_37[171]    = ( l_38 [324] & !i[1815]) | ( l_38 [325] &  i[1815]);
assign l_37[172]    = ( l_38 [326] & !i[1815]) | ( l_38 [327] &  i[1815]);
assign l_37[173]    = ( l_38 [328] & !i[1815]) | ( l_38 [329] &  i[1815]);
assign l_37[174]    = ( l_38 [330] & !i[1815]) | ( l_38 [331] &  i[1815]);
assign l_37[175]    = ( l_38 [332] & !i[1815]) | ( l_38 [333] &  i[1815]);
assign l_37[176]    = ( l_38 [334] & !i[1815]) | ( l_38 [335] &  i[1815]);
assign l_37[177]    = ( l_38 [336] & !i[1815]) | ( l_38 [337] &  i[1815]);
assign l_37[178]    = ( l_38 [338] & !i[1815]) | ( l_38 [339] &  i[1815]);
assign l_37[179]    = ( l_38 [340] & !i[1815]) | ( l_38 [341] &  i[1815]);
assign l_37[180]    = ( l_38 [342] & !i[1815]) | ( l_38 [343] &  i[1815]);
assign l_37[181]    = ( l_38 [344] & !i[1815]) | ( l_38 [345] &  i[1815]);
assign l_37[182]    = ( l_38 [346] & !i[1815]) | ( l_38 [347] &  i[1815]);
assign l_37[183]    = ( l_38 [348] & !i[1815]) | ( l_38 [349] &  i[1815]);
assign l_37[184]    = ( l_38 [350] & !i[1815]) | ( l_38 [351] &  i[1815]);
assign l_37[185]    = ( l_38 [352] & !i[1815]) | ( l_38 [353] &  i[1815]);
assign l_37[186]    = ( l_38 [354] & !i[1815]) | ( l_38 [355] &  i[1815]);
assign l_37[187]    = ( l_38 [356] & !i[1815]) | ( l_38 [357] &  i[1815]);
assign l_37[188]    = ( l_38 [358] & !i[1815]) | ( l_38 [359] &  i[1815]);
assign l_37[189]    = ( l_38 [360] & !i[1815]) | ( l_38 [361] &  i[1815]);
assign l_37[190]    = ( l_38 [362] & !i[1815]) | ( l_38 [363] &  i[1815]);
assign l_37[191]    = ( l_38 [364] & !i[1815]) | ( l_38 [365] &  i[1815]);
assign l_37[192]    = ( l_38 [366] & !i[1815]) | ( l_38 [367] &  i[1815]);
assign l_37[193]    = ( l_38 [368] & !i[1815]) | ( l_38 [369] &  i[1815]);
assign l_37[194]    = ( l_38 [370] & !i[1815]) | ( l_38 [371] &  i[1815]);
assign l_37[195]    = ( l_38 [372] & !i[1815]) | ( l_38 [373] &  i[1815]);
assign l_37[196]    = ( l_38 [374] & !i[1815]) | ( l_38 [375] &  i[1815]);
assign l_37[197]    = ( l_38 [376] & !i[1815]) | ( l_38 [377] &  i[1815]);
assign l_37[198]    = ( l_38 [378] & !i[1815]) | ( l_38 [379] &  i[1815]);
assign l_37[199]    = ( l_38 [380] & !i[1815]) | ( l_38 [381] &  i[1815]);
assign l_37[200]    = ( l_38 [382] & !i[1815]) | ( l_38 [383] &  i[1815]);
assign l_37[201]    = ( l_38 [384] & !i[1815]) | ( l_38 [385] &  i[1815]);
assign l_37[202]    = ( l_38 [386] & !i[1815]) | ( l_38 [387] &  i[1815]);
assign l_37[203]    = ( l_38 [388] & !i[1815]) | ( l_38 [389] &  i[1815]);
assign l_37[204]    = ( l_38 [390] & !i[1815]) | ( l_38 [391] &  i[1815]);
assign l_37[205]    = ( l_38 [392] & !i[1815]) | ( l_38 [393] &  i[1815]);
assign l_37[206]    = ( l_38 [394] & !i[1815]) | ( l_38 [395] &  i[1815]);
assign l_37[207]    = ( l_38 [396] & !i[1815]) | ( l_38 [397] &  i[1815]);
assign l_37[208]    = ( l_38 [398] & !i[1815]) | ( l_38 [399] &  i[1815]);
assign l_37[209]    = ( l_38 [400] & !i[1815]) | ( l_38 [401] &  i[1815]);
assign l_37[210]    = ( l_38 [402] & !i[1815]) | ( l_38 [403] &  i[1815]);
assign l_37[211]    = ( l_38 [404] & !i[1815]) | ( l_38 [405] &  i[1815]);
assign l_37[212]    = ( l_38 [406] & !i[1815]) | ( l_38 [407] &  i[1815]);
assign l_37[213]    = ( l_38 [408] & !i[1815]) | ( l_38 [409] &  i[1815]);
assign l_37[214]    = ( l_38 [410] & !i[1815]) | ( l_38 [411] &  i[1815]);
assign l_37[215]    = ( l_38 [412] & !i[1815]) | ( l_38 [413] &  i[1815]);
assign l_37[216]    = ( l_38 [414] & !i[1815]) | ( l_38 [415] &  i[1815]);
assign l_37[217]    = ( l_38 [416] & !i[1815]) | ( l_38 [417] &  i[1815]);
assign l_37[218]    = ( l_38 [418] & !i[1815]) | ( l_38 [419] &  i[1815]);
assign l_37[219]    = ( l_38 [420] & !i[1815]) | ( l_38 [421] &  i[1815]);
assign l_37[220]    = ( l_38 [422] & !i[1815]) | ( l_38 [423] &  i[1815]);
assign l_37[221]    = ( l_38 [424] & !i[1815]) | ( l_38 [425] &  i[1815]);
assign l_37[222]    = ( l_38 [426] & !i[1815]) | ( l_38 [427] &  i[1815]);
assign l_37[223]    = ( l_38 [428] & !i[1815]) | ( l_38 [429] &  i[1815]);
assign l_37[224]    = ( l_38 [430] & !i[1815]) | ( l_38 [431] &  i[1815]);
assign l_37[225]    = ( l_38 [432] & !i[1815]) | ( l_38 [433] &  i[1815]);
assign l_37[226]    = ( l_38 [434] & !i[1815]) | ( l_38 [435] &  i[1815]);
assign l_37[227]    = ( l_38 [436] & !i[1815]) | ( l_38 [437] &  i[1815]);
assign l_37[228]    = ( l_38 [438] & !i[1815]) | ( l_38 [439] &  i[1815]);
assign l_37[229]    = ( l_38 [440] & !i[1815]) | ( l_38 [441] &  i[1815]);
assign l_37[230]    = ( l_38 [442] & !i[1815]) | ( l_38 [443] &  i[1815]);
assign l_37[231]    = ( l_38 [444] & !i[1815]) | ( l_38 [445] &  i[1815]);
assign l_37[232]    = ( l_38 [446] & !i[1815]) | ( l_38 [447] &  i[1815]);
assign l_37[233]    = ( l_38 [448] & !i[1815]) | ( l_38 [449] &  i[1815]);
assign l_37[234]    = ( l_38 [450] & !i[1815]) | ( l_38 [451] &  i[1815]);
assign l_37[235]    = ( l_38 [452] & !i[1815]) | ( l_38 [453] &  i[1815]);
assign l_37[236]    = ( l_38 [454] & !i[1815]) | ( l_38 [455] &  i[1815]);
assign l_37[237]    = ( l_38 [456] & !i[1815]) | ( l_38 [457] &  i[1815]);
assign l_37[238]    = ( l_38 [458] & !i[1815]) | ( l_38 [459] &  i[1815]);
assign l_37[239]    = ( l_38 [460] & !i[1815]) | ( l_38 [461] &  i[1815]);
assign l_37[240]    = ( l_38 [462] & !i[1815]) | ( l_38 [463] &  i[1815]);
assign l_37[241]    = ( l_38 [464] & !i[1815]) | ( l_38 [465] &  i[1815]);
assign l_37[242]    = ( l_38 [466] & !i[1815]) | ( l_38 [467] &  i[1815]);
assign l_37[243]    = ( l_38 [468] & !i[1815]) | ( l_38 [469] &  i[1815]);
assign l_37[244]    = ( l_38 [470] & !i[1815]) | ( l_38 [471] &  i[1815]);
assign l_37[245]    = ( l_38 [472] & !i[1815]) | ( l_38 [473] &  i[1815]);
assign l_37[246]    = ( l_38 [474] & !i[1815]) | ( l_38 [475] &  i[1815]);
assign l_37[247]    = ( l_38 [476] & !i[1815]) | ( l_38 [477] &  i[1815]);
assign l_37[248]    = ( l_38 [478] & !i[1815]) | ( l_38 [479] &  i[1815]);
assign l_37[249]    = ( l_38 [480] & !i[1815]) | ( l_38 [481] &  i[1815]);
assign l_37[250]    = ( l_38 [482] & !i[1815]) | ( l_38 [483] &  i[1815]);
assign l_37[251]    = ( l_38 [484] & !i[1815]) | ( l_38 [485] &  i[1815]);
assign l_37[252]    = ( l_38 [486] & !i[1815]) | ( l_38 [487] &  i[1815]);
assign l_37[253]    = ( l_38 [488] & !i[1815]) | ( l_38 [489] &  i[1815]);
assign l_37[254]    = ( l_38 [490] & !i[1815]) | ( l_38 [491] &  i[1815]);
assign l_37[255]    = ( l_38 [492] & !i[1815]) | ( l_38 [493] &  i[1815]);
assign l_37[256]    = ( l_38 [494] & !i[1815]) | ( l_38 [495] &  i[1815]);
assign l_37[257]    = ( l_38 [496] & !i[1815]) | ( l_38 [497] &  i[1815]);
assign l_37[258]    = ( l_38 [498] & !i[1815]) | ( l_38 [499] &  i[1815]);
assign l_37[259]    = ( l_38 [500] & !i[1815]) | ( l_38 [501] &  i[1815]);
assign l_37[260]    = ( l_38 [502] & !i[1815]) | ( l_38 [503] &  i[1815]);
assign l_37[261]    = ( l_38 [504] & !i[1815]) | ( l_38 [505] &  i[1815]);
assign l_37[262]    = ( l_38 [506] & !i[1815]) | ( l_38 [507] &  i[1815]);
assign l_37[263]    = ( l_38 [508] & !i[1815]) | ( l_38 [509] &  i[1815]);
assign l_37[264]    = ( l_38 [510] & !i[1815]) | ( l_38 [511] &  i[1815]);
assign l_37[265]    = ( l_38 [512] & !i[1815]) | ( l_38 [513] &  i[1815]);
assign l_37[266]    = ( l_38 [514] & !i[1815]) | ( l_38 [515] &  i[1815]);
assign l_37[267]    = ( l_38 [516] & !i[1815]) | ( l_38 [517] &  i[1815]);
assign l_37[268]    = ( l_38 [518] & !i[1815]) | ( l_38 [519] &  i[1815]);
assign l_37[269]    = ( l_38 [520] & !i[1815]) | ( l_38 [521] &  i[1815]);
assign l_37[270]    = ( l_38 [522] & !i[1815]) | ( l_38 [523] &  i[1815]);
assign l_37[271]    = ( l_38 [524] & !i[1815]) | ( l_38 [525] &  i[1815]);
assign l_37[272]    = ( l_38 [526] & !i[1815]) | ( l_38 [527] &  i[1815]);
assign l_37[273]    = ( l_38 [528] & !i[1815]) | ( l_38 [529] &  i[1815]);
assign l_37[274]    = ( l_38 [530] & !i[1815]) | ( l_38 [531] &  i[1815]);
assign l_37[275]    = ( l_38 [532] & !i[1815]) | ( l_38 [533] &  i[1815]);
assign l_37[276]    = ( l_38 [534] & !i[1815]) | ( l_38 [535] &  i[1815]);
assign l_37[277]    = ( l_38 [536] & !i[1815]) | ( l_38 [537] &  i[1815]);
assign l_37[278]    = ( l_38 [538] & !i[1815]) | ( l_38 [539] &  i[1815]);
assign l_37[279]    = ( l_38 [540] & !i[1815]) | ( l_38 [541] &  i[1815]);
assign l_37[280]    = ( l_38 [542] & !i[1815]) | ( l_38 [543] &  i[1815]);
assign l_37[281]    = ( l_38 [544] & !i[1815]) | ( l_38 [545] &  i[1815]);
assign l_37[282]    = ( l_38 [546] & !i[1815]) | ( l_38 [547] &  i[1815]);
assign l_37[283]    = ( l_38 [548] & !i[1815]) | ( l_38 [549] &  i[1815]);
assign l_37[284]    = ( l_38 [550] & !i[1815]) | ( l_38 [551] &  i[1815]);
assign l_37[285]    = ( l_38 [552] & !i[1815]) | ( l_38 [553] &  i[1815]);
assign l_37[286]    = ( l_38 [554] & !i[1815]) | ( l_38 [555] &  i[1815]);
assign l_37[287]    = ( l_38 [556] & !i[1815]) | ( l_38 [557] &  i[1815]);
assign l_37[288]    = ( l_38 [558] & !i[1815]) | ( l_38 [559] &  i[1815]);
assign l_37[289]    = ( l_38 [560] & !i[1815]) | ( l_38 [561] &  i[1815]);
assign l_37[290]    = ( l_38 [562] & !i[1815]) | ( l_38 [563] &  i[1815]);
assign l_37[291]    = ( l_38 [564] & !i[1815]) | ( l_38 [565] &  i[1815]);
assign l_37[292]    = ( l_38 [566] & !i[1815]) | ( l_38 [567] &  i[1815]);
assign l_37[293]    = ( l_38 [568] & !i[1815]) | ( l_38 [569] &  i[1815]);
assign l_37[294]    = ( l_38 [570] & !i[1815]) | ( l_38 [571] &  i[1815]);
assign l_37[295]    = ( l_38 [572] & !i[1815]) | ( l_38 [573] &  i[1815]);
assign l_37[296]    = ( l_38 [574] & !i[1815]) | ( l_38 [575] &  i[1815]);
assign l_37[297]    = ( l_38 [576] & !i[1815]) | ( l_38 [577] &  i[1815]);
assign l_37[298]    = ( l_38 [578] & !i[1815]) | ( l_38 [579] &  i[1815]);
assign l_37[299]    = ( l_38 [580] & !i[1815]) | ( l_38 [581] &  i[1815]);
assign l_37[300]    = ( l_38 [582] & !i[1815]) | ( l_38 [583] &  i[1815]);
assign l_37[301]    = ( l_38 [584] & !i[1815]) | ( l_38 [585] &  i[1815]);
assign l_37[302]    = ( l_38 [586] & !i[1815]) | ( l_38 [587] &  i[1815]);
assign l_37[303]    = ( l_38 [588] & !i[1815]) | ( l_38 [589] &  i[1815]);
assign l_37[304]    = ( l_38 [590] & !i[1815]) | ( l_38 [591] &  i[1815]);
assign l_37[305]    = ( l_38 [592] & !i[1815]) | ( l_38 [593] &  i[1815]);
assign l_37[306]    = ( l_38 [594] & !i[1815]) | ( l_38 [595] &  i[1815]);
assign l_37[307]    = ( l_38 [596] & !i[1815]) | ( l_38 [597] &  i[1815]);
assign l_37[308]    = ( l_38 [598] & !i[1815]) | ( l_38 [599] &  i[1815]);
assign l_37[309]    = ( l_38 [600] & !i[1815]) | ( l_38 [601] &  i[1815]);
assign l_37[310]    = ( l_38 [602] & !i[1815]) | ( l_38 [603] &  i[1815]);
assign l_37[311]    = ( l_38 [604] & !i[1815]) | ( l_38 [605] &  i[1815]);
assign l_37[312]    = ( l_38 [606] & !i[1815]) | ( l_38 [607] &  i[1815]);
assign l_37[313]    = ( l_38 [608] & !i[1815]) | ( l_38 [609] &  i[1815]);
assign l_37[314]    = ( l_38 [610] & !i[1815]) | ( l_38 [611] &  i[1815]);
assign l_37[315]    = ( l_38 [612] & !i[1815]) | ( l_38 [613] &  i[1815]);
assign l_37[316]    = ( l_38 [614] & !i[1815]) | ( l_38 [615] &  i[1815]);
assign l_37[317]    = ( l_38 [616] & !i[1815]) | ( l_38 [617] &  i[1815]);
assign l_37[318]    = ( l_38 [618] & !i[1815]) | ( l_38 [619] &  i[1815]);
assign l_37[319]    = ( l_38 [620] & !i[1815]) | ( l_38 [621] &  i[1815]);
assign l_37[320]    = ( l_38 [622] & !i[1815]) | ( l_38 [623] &  i[1815]);
assign l_37[321]    = ( l_38 [624] & !i[1815]) | ( l_38 [625] &  i[1815]);
assign l_37[322]    = ( l_38 [626] & !i[1815]) | ( l_38 [627] &  i[1815]);
assign l_37[323]    = ( l_38 [628] & !i[1815]) | ( l_38 [629] &  i[1815]);
assign l_37[324]    = ( l_38 [630] & !i[1815]) | ( l_38 [631] &  i[1815]);
assign l_37[325]    = ( l_38 [632] & !i[1815]) | ( l_38 [633] &  i[1815]);
assign l_37[326]    = ( l_38 [634] & !i[1815]) | ( l_38 [635] &  i[1815]);
assign l_37[327]    = ( l_38 [636] & !i[1815]) | ( l_38 [637] &  i[1815]);
assign l_37[328]    = ( l_38 [638] & !i[1815]) | ( l_38 [639] &  i[1815]);
assign l_37[329]    = ( l_38 [640] & !i[1815]) | ( l_38 [641] &  i[1815]);
assign l_37[330]    = ( l_38 [642] & !i[1815]) | ( l_38 [643] &  i[1815]);
assign l_37[331]    = ( l_38 [644] & !i[1815]) | ( l_38 [645] &  i[1815]);
assign l_37[332]    = ( l_38 [646] & !i[1815]) | ( l_38 [647] &  i[1815]);
assign l_37[333]    = ( l_38 [648] & !i[1815]) | ( l_38 [649] &  i[1815]);
assign l_37[334]    = ( l_38 [650] & !i[1815]) | ( l_38 [651] &  i[1815]);
assign l_37[335]    = ( l_38 [652] & !i[1815]) | ( l_38 [653] &  i[1815]);
assign l_37[336]    = ( l_38 [654] & !i[1815]) | ( l_38 [655] &  i[1815]);
assign l_37[337]    = ( l_38 [656] & !i[1815]) | ( l_38 [657] &  i[1815]);
assign l_37[338]    = ( l_38 [658] & !i[1815]) | ( l_38 [659] &  i[1815]);
assign l_37[339]    = ( l_38 [660] & !i[1815]) | ( l_38 [661] &  i[1815]);
assign l_37[340]    = ( l_38 [662] & !i[1815]) | ( l_38 [663] &  i[1815]);
assign l_37[341]    = ( l_38 [664] & !i[1815]) | ( l_38 [665] &  i[1815]);
assign l_37[342]    = ( l_38 [666] & !i[1815]) | ( l_38 [667] &  i[1815]);
assign l_37[343]    = ( l_38 [668] & !i[1815]) | ( l_38 [669] &  i[1815]);
assign l_37[344]    = ( l_38 [670] & !i[1815]) | ( l_38 [671] &  i[1815]);
assign l_37[345]    = ( l_38 [672] & !i[1815]) | ( l_38 [673] &  i[1815]);
assign l_37[346]    = ( l_38 [674] & !i[1815]) | ( l_38 [675] &  i[1815]);
assign l_37[347]    = ( l_38 [676] & !i[1815]) | ( l_38 [677] &  i[1815]);
assign l_37[348]    = ( l_38 [678] & !i[1815]) | ( l_38 [679] &  i[1815]);
assign l_37[349]    = ( l_38 [680] & !i[1815]) | ( l_38 [681] &  i[1815]);
assign l_37[350]    = ( l_38 [682] & !i[1815]) | ( l_38 [683] &  i[1815]);
assign l_37[351]    = ( l_38 [684] & !i[1815]) | ( l_38 [685] &  i[1815]);
assign l_37[352]    = ( l_38 [686] & !i[1815]) | ( l_38 [687] &  i[1815]);
assign l_37[353]    = ( l_38 [688] & !i[1815]) | ( l_38 [689] &  i[1815]);
assign l_37[354]    = ( l_38 [690] & !i[1815]) | ( l_38 [691] &  i[1815]);
assign l_37[355]    = ( l_38 [692] & !i[1815]) | ( l_38 [693] &  i[1815]);
assign l_37[356]    = ( l_38 [694] & !i[1815]) | ( l_38 [695] &  i[1815]);
assign l_37[357]    = ( l_38 [696] & !i[1815]) | ( l_38 [697] &  i[1815]);
assign l_37[358]    = ( l_38 [698] & !i[1815]) | ( l_38 [699] &  i[1815]);
assign l_37[359]    = ( l_38 [700] & !i[1815]) | ( l_38 [701] &  i[1815]);
assign l_37[360]    = ( l_38 [702] & !i[1815]) | ( l_38 [703] &  i[1815]);
assign l_37[361]    = ( l_38 [704] & !i[1815]) | ( l_38 [705] &  i[1815]);
assign l_37[362]    = ( l_38 [706] & !i[1815]) | ( l_38 [707] &  i[1815]);
assign l_37[363]    = ( l_38 [708] & !i[1815]) | ( l_38 [709] &  i[1815]);
assign l_37[364]    = ( l_38 [710] & !i[1815]) | ( l_38 [711] &  i[1815]);
assign l_37[365]    = ( l_38 [712] & !i[1815]) | ( l_38 [713] &  i[1815]);
assign l_37[366]    = ( l_38 [714] & !i[1815]) | ( l_38 [715] &  i[1815]);
assign l_37[367]    = ( l_38 [716] & !i[1815]) | ( l_38 [717] &  i[1815]);
assign l_37[368]    = ( l_38 [718] & !i[1815]) | ( l_38 [719] &  i[1815]);
assign l_37[369]    = ( l_38 [720] & !i[1815]) | ( l_38 [721] &  i[1815]);
assign l_37[370]    = ( l_38 [722] & !i[1815]) | ( l_38 [723] &  i[1815]);
assign l_37[371]    = ( l_38 [724] & !i[1815]) | ( l_38 [725] &  i[1815]);
assign l_37[372]    = ( l_38 [726] & !i[1815]) | ( l_38 [727] &  i[1815]);
assign l_37[373]    = ( l_38 [728] & !i[1815]) | ( l_38 [729] &  i[1815]);
assign l_37[374]    = ( l_38 [730] & !i[1815]) | ( l_38 [731] &  i[1815]);
assign l_37[375]    = ( l_38 [732] & !i[1815]) | ( l_38 [733] &  i[1815]);
assign l_37[376]    = ( l_38 [734] & !i[1815]) | ( l_38 [735] &  i[1815]);
assign l_37[377]    = ( l_38 [736] & !i[1815]) | ( l_38 [737] &  i[1815]);
assign l_37[378]    = ( l_38 [738] & !i[1815]) | ( l_38 [739] &  i[1815]);
assign l_37[379]    = ( l_38 [740] & !i[1815]) | ( l_38 [741] &  i[1815]);
assign l_37[380]    = ( l_38 [742] & !i[1815]) | ( l_38 [743] &  i[1815]);
assign l_37[381]    = ( l_38 [744] & !i[1815]) | ( l_38 [745] &  i[1815]);
assign l_37[382]    = ( l_38 [746] & !i[1815]) | ( l_38 [747] &  i[1815]);
assign l_37[383]    = ( l_38 [748] & !i[1815]) | ( l_38 [749] &  i[1815]);
assign l_37[384]    = ( l_38 [750] & !i[1815]) | ( l_38 [751] &  i[1815]);
assign l_37[385]    = ( l_38 [752] & !i[1815]) | ( l_38 [753] &  i[1815]);
assign l_37[386]    = ( l_38 [754] & !i[1815]) | ( l_38 [755] &  i[1815]);
assign l_37[387]    = ( l_38 [756] & !i[1815]) | ( l_38 [757] &  i[1815]);
assign l_37[388]    = ( l_38 [758] & !i[1815]) | ( l_38 [759] &  i[1815]);
assign l_37[389]    = ( l_38 [760] & !i[1815]) | ( l_38 [761] &  i[1815]);
assign l_37[390]    = ( l_38 [762] & !i[1815]) | ( l_38 [763] &  i[1815]);
assign l_37[391]    = ( l_38 [764] & !i[1815]) | ( l_38 [765] &  i[1815]);
assign l_37[392]    = ( l_38 [766] & !i[1815]) | ( l_38 [767] &  i[1815]);
assign l_37[393]    = ( l_38 [768] & !i[1815]) | ( l_38 [769] &  i[1815]);
assign l_37[394]    = ( l_38 [770] & !i[1815]) | ( l_38 [771] &  i[1815]);
assign l_37[395]    = ( l_38 [772] & !i[1815]) | ( l_38 [773] &  i[1815]);
assign l_37[396]    = ( l_38 [774] & !i[1815]) | ( l_38 [775] &  i[1815]);
assign l_37[397]    = ( l_38 [776] & !i[1815]) | ( l_38 [777] &  i[1815]);
assign l_37[398]    = ( l_38 [778] & !i[1815]) | ( l_38 [779] &  i[1815]);
assign l_37[399]    = ( l_38 [780] & !i[1815]) | ( l_38 [781] &  i[1815]);
assign l_37[400]    = ( l_38 [782] & !i[1815]) | ( l_38 [783] &  i[1815]);
assign l_37[401]    = ( l_38 [784] & !i[1815]) | ( l_38 [785] &  i[1815]);
assign l_37[402]    = ( l_38 [786] & !i[1815]) | ( l_38 [787] &  i[1815]);
assign l_37[403]    = ( l_38 [788] & !i[1815]) | ( l_38 [789] &  i[1815]);
assign l_37[404]    = ( l_38 [790] & !i[1815]) | ( l_38 [791] &  i[1815]);
assign l_37[405]    = ( l_38 [792] & !i[1815]) | ( l_38 [793] &  i[1815]);
assign l_37[406]    = ( l_38 [794] & !i[1815]) | ( l_38 [795] &  i[1815]);
assign l_37[407]    = ( l_38 [796] & !i[1815]) | ( l_38 [797] &  i[1815]);
assign l_37[408]    = ( l_38 [798] & !i[1815]) | ( l_38 [799] &  i[1815]);
assign l_37[409]    = ( l_38 [800] & !i[1815]) | ( l_38 [801] &  i[1815]);
assign l_37[410]    = ( l_38 [802] & !i[1815]) | ( l_38 [803] &  i[1815]);
assign l_37[411]    = ( l_38 [804] & !i[1815]) | ( l_38 [805] &  i[1815]);
assign l_37[412]    = ( l_38 [806] & !i[1815]) | ( l_38 [807] &  i[1815]);
assign l_37[413]    = ( l_38 [808] & !i[1815]) | ( l_38 [809] &  i[1815]);
assign l_37[414]    = ( l_38 [810] & !i[1815]) | ( l_38 [811] &  i[1815]);
assign l_37[415]    = ( l_38 [812] & !i[1815]) | ( l_38 [813] &  i[1815]);
assign l_37[416]    = ( l_38 [814] & !i[1815]) | ( l_38 [815] &  i[1815]);
assign l_37[417]    = ( l_38 [816] & !i[1815]) | ( l_38 [817] &  i[1815]);
assign l_37[418]    = ( l_38 [818] & !i[1815]) | ( l_38 [819] &  i[1815]);
assign l_37[419]    = ( l_38 [820] & !i[1815]) | ( l_38 [821] &  i[1815]);
assign l_37[420]    = ( l_38 [822] & !i[1815]) | ( l_38 [823] &  i[1815]);
assign l_37[421]    = ( l_38 [824] & !i[1815]) | ( l_38 [825] &  i[1815]);
assign l_37[422]    = ( l_38 [826] & !i[1815]) | ( l_38 [827] &  i[1815]);
assign l_37[423]    = ( l_38 [828] & !i[1815]) | ( l_38 [829] &  i[1815]);
assign l_37[424]    = ( l_38 [830] & !i[1815]) | ( l_38 [831] &  i[1815]);
assign l_37[425]    = ( l_38 [832] & !i[1815]) | ( l_38 [833] &  i[1815]);
assign l_37[426]    = ( l_38 [834] & !i[1815]) | ( l_38 [835] &  i[1815]);
assign l_37[427]    = ( l_38 [836] & !i[1815]) | ( l_38 [837] &  i[1815]);
assign l_37[428]    = ( l_38 [838] & !i[1815]) | ( l_38 [839] &  i[1815]);
assign l_37[429]    = ( l_38 [840] & !i[1815]) | ( l_38 [841] &  i[1815]);
assign l_37[430]    = ( l_38 [842] & !i[1815]) | ( l_38 [843] &  i[1815]);
assign l_37[431]    = ( l_38 [844] & !i[1815]) | ( l_38 [845] &  i[1815]);
assign l_37[432]    = ( l_38 [846] & !i[1815]) | ( l_38 [847] &  i[1815]);
assign l_37[433]    = ( l_38 [848] & !i[1815]) | ( l_38 [849] &  i[1815]);
assign l_37[434]    = ( l_38 [850] & !i[1815]) | ( l_38 [851] &  i[1815]);
assign l_37[435]    = ( l_38 [852] & !i[1815]) | ( l_38 [853] &  i[1815]);
assign l_37[436]    = ( l_38 [854] & !i[1815]) | ( l_38 [855] &  i[1815]);
assign l_37[437]    = ( l_38 [856] & !i[1815]) | ( l_38 [857] &  i[1815]);
assign l_37[438]    = ( l_38 [858] & !i[1815]) | ( l_38 [859] &  i[1815]);
assign l_37[439]    = ( l_38 [860] & !i[1815]) | ( l_38 [861] &  i[1815]);
assign l_37[440]    = ( l_38 [862] & !i[1815]) | ( l_38 [863] &  i[1815]);
assign l_37[441]    = ( l_38 [864] & !i[1815]) | ( l_38 [865] &  i[1815]);
assign l_37[442]    = ( l_38 [866] & !i[1815]) | ( l_38 [867] &  i[1815]);
assign l_37[443]    = ( l_38 [868] & !i[1815]) | ( l_38 [869] &  i[1815]);
assign l_37[444]    = ( l_38 [870] & !i[1815]) | ( l_38 [871] &  i[1815]);
assign l_37[445]    = ( l_38 [872] & !i[1815]) | ( l_38 [873] &  i[1815]);
assign l_37[446]    = ( l_38 [874] & !i[1815]) | ( l_38 [875] &  i[1815]);
assign l_37[447]    = ( l_38 [876] & !i[1815]) | ( l_38 [877] &  i[1815]);
assign l_37[448]    = ( l_38 [878] & !i[1815]) | ( l_38 [879] &  i[1815]);
assign l_37[449]    = ( l_38 [880] & !i[1815]) | ( l_38 [881] &  i[1815]);
assign l_37[450]    = ( l_38 [882] & !i[1815]) | ( l_38 [883] &  i[1815]);
assign l_37[451]    = ( l_38 [884] & !i[1815]) | ( l_38 [885] &  i[1815]);
assign l_37[452]    = ( l_38 [886] & !i[1815]) | ( l_38 [887] &  i[1815]);
assign l_37[453]    = ( l_38 [888] & !i[1815]) | ( l_38 [889] &  i[1815]);
assign l_37[454]    = ( l_38 [890] & !i[1815]) | ( l_38 [891] &  i[1815]);
assign l_37[455]    = ( l_38 [892] & !i[1815]) | ( l_38 [893] &  i[1815]);
assign l_37[456]    = ( l_38 [894] & !i[1815]) | ( l_38 [895] &  i[1815]);
assign l_37[457]    = ( l_38 [896] & !i[1815]) | ( l_38 [897] &  i[1815]);
assign l_37[458]    = ( l_38 [898] & !i[1815]) | ( l_38 [899] &  i[1815]);
assign l_37[459]    = ( l_38 [900] & !i[1815]) | ( l_38 [901] &  i[1815]);
assign l_37[460]    = ( l_38 [902] & !i[1815]) | ( l_38 [903] &  i[1815]);
assign l_37[461]    = ( l_38 [904] & !i[1815]) | ( l_38 [905] &  i[1815]);
assign l_37[462]    = ( l_38 [906] & !i[1815]) | ( l_38 [907] &  i[1815]);
assign l_37[463]    = ( l_38 [908] & !i[1815]) | ( l_38 [909] &  i[1815]);
assign l_37[464]    = ( l_38 [910] & !i[1815]) | ( l_38 [911] &  i[1815]);
assign l_37[465]    = ( l_38 [912] & !i[1815]) | ( l_38 [913] &  i[1815]);
assign l_37[466]    = ( l_38 [914] & !i[1815]) | ( l_38 [915] &  i[1815]);
assign l_37[467]    = ( l_38 [916] & !i[1815]) | ( l_38 [917] &  i[1815]);
assign l_37[468]    = ( l_38 [918] & !i[1815]) | ( l_38 [919] &  i[1815]);
assign l_37[469]    = ( l_38 [920] & !i[1815]) | ( l_38 [921] &  i[1815]);
assign l_37[470]    = ( l_38 [922] & !i[1815]) | ( l_38 [923] &  i[1815]);
assign l_37[471]    = ( l_38 [924] & !i[1815]) | ( l_38 [925] &  i[1815]);
assign l_37[472]    = ( l_38 [926] & !i[1815]) | ( l_38 [927] &  i[1815]);
assign l_37[473]    = ( l_38 [928] & !i[1815]) | ( l_38 [929] &  i[1815]);
assign l_37[474]    = ( l_38 [930] & !i[1815]) | ( l_38 [931] &  i[1815]);
assign l_37[475]    = ( l_38 [932] & !i[1815]) | ( l_38 [933] &  i[1815]);
assign l_37[476]    = ( l_38 [934] & !i[1815]) | ( l_38 [935] &  i[1815]);
assign l_37[477]    = ( l_38 [936] & !i[1815]) | ( l_38 [937] &  i[1815]);
assign l_37[478]    = ( l_38 [938] & !i[1815]) | ( l_38 [939] &  i[1815]);
assign l_37[479]    = ( l_38 [940] & !i[1815]) | ( l_38 [941] &  i[1815]);
assign l_37[480]    = ( l_38 [942] & !i[1815]) | ( l_38 [943] &  i[1815]);
assign l_37[481]    = ( l_38 [944] & !i[1815]) | ( l_38 [945] &  i[1815]);
assign l_37[482]    = ( l_38 [946] & !i[1815]) | ( l_38 [947] &  i[1815]);
assign l_37[483]    = ( l_38 [948] & !i[1815]) | ( l_38 [949] &  i[1815]);
assign l_37[484]    = ( l_38 [950] & !i[1815]) | ( l_38 [951] &  i[1815]);
assign l_37[485]    = ( l_38 [952] & !i[1815]) | ( l_38 [953] &  i[1815]);
assign l_37[486]    = ( l_38 [954] & !i[1815]) | ( l_38 [955] &  i[1815]);
assign l_37[487]    = ( l_38 [956] & !i[1815]) | ( l_38 [957] &  i[1815]);
assign l_37[488]    = ( l_38 [958] & !i[1815]) | ( l_38 [959] &  i[1815]);
assign l_37[489]    = ( l_38 [960] & !i[1815]) | ( l_38 [961] &  i[1815]);
assign l_37[490]    = ( l_38 [962] & !i[1815]) | ( l_38 [963] &  i[1815]);
assign l_37[491]    = ( l_38 [964] & !i[1815]) | ( l_38 [965] &  i[1815]);
assign l_37[492]    = ( l_38 [966] & !i[1815]) | ( l_38 [967] &  i[1815]);
assign l_37[493]    = ( l_38 [968] & !i[1815]) | ( l_38 [969] &  i[1815]);
assign l_37[494]    = ( l_38 [970] & !i[1815]) | ( l_38 [971] &  i[1815]);
assign l_37[495]    = ( l_38 [972] & !i[1815]) | ( l_38 [973] &  i[1815]);
assign l_37[496]    = ( l_38 [974] & !i[1815]) | ( l_38 [975] &  i[1815]);
assign l_37[497]    = ( l_38 [976] & !i[1815]) | ( l_38 [977] &  i[1815]);
assign l_37[498]    = ( l_38 [978] & !i[1815]) | ( l_38 [979] &  i[1815]);
assign l_37[499]    = ( l_38 [980] & !i[1815]) | ( l_38 [981] &  i[1815]);
assign l_37[500]    = ( l_38 [982] & !i[1815]) | ( l_38 [983] &  i[1815]);
assign l_37[501]    = ( l_38 [984] & !i[1815]) | ( l_38 [985] &  i[1815]);
assign l_37[502]    = ( l_38 [986] & !i[1815]) | ( l_38 [987] &  i[1815]);
assign l_37[503]    = ( l_38 [988] & !i[1815]) | ( l_38 [989] &  i[1815]);
assign l_37[504]    = ( l_38 [990] & !i[1815]) | ( l_38 [991] &  i[1815]);
assign l_37[505]    = ( l_38 [992] & !i[1815]) | ( l_38 [993] &  i[1815]);
assign l_37[506]    = ( l_38 [994] & !i[1815]) | ( l_38 [995] &  i[1815]);
assign l_37[507]    = ( l_38 [996] & !i[1815]) | ( l_38 [997] &  i[1815]);
assign l_37[508]    = ( l_38 [998] & !i[1815]) | ( l_38 [999] &  i[1815]);
assign l_37[509]    = ( l_38 [1000] & !i[1815]) | ( l_38 [1001] &  i[1815]);
assign l_37[510]    = ( l_38 [1002] & !i[1815]) | ( l_38 [1003] &  i[1815]);
assign l_37[511]    = ( l_38 [1004] & !i[1815]) | ( l_38 [1005] &  i[1815]);
assign l_37[512]    = ( l_38 [1006] & !i[1815]) | ( l_38 [1007] &  i[1815]);
assign l_37[513]    = ( l_38 [1008] & !i[1815]) | ( l_38 [1009] &  i[1815]);
assign l_37[514]    = ( l_38 [1010] & !i[1815]) | ( l_38 [1011] &  i[1815]);
assign l_37[515]    = ( l_38 [1012] & !i[1815]) | ( l_38 [1013] &  i[1815]);
assign l_37[516]    = ( l_38 [1014] & !i[1815]) | ( l_38 [1015] &  i[1815]);
assign l_37[517]    = ( l_38 [1016] & !i[1815]) | ( l_38 [1017] &  i[1815]);
assign l_37[518]    = ( l_38 [1018] & !i[1815]) | ( l_38 [1019] &  i[1815]);
assign l_37[519]    = ( l_38 [1020] & !i[1815]) | ( l_38 [1021] &  i[1815]);
assign l_37[520]    = ( l_38 [1022] & !i[1815]) | ( l_38 [1023] &  i[1815]);
assign l_37[521]    = ( l_38 [1024] & !i[1815]) | ( l_38 [1025] &  i[1815]);
assign l_37[522]    = ( l_38 [1026] & !i[1815]) | ( l_38 [1027] &  i[1815]);
assign l_37[523]    = ( l_38 [1028] & !i[1815]) | ( l_38 [1029] &  i[1815]);
assign l_37[524]    = ( l_38 [1030] & !i[1815]) | ( l_38 [1031] &  i[1815]);
assign l_37[525]    = ( l_38 [1032] & !i[1815]) | ( l_38 [1033] &  i[1815]);
assign l_37[526]    = ( l_38 [1034] & !i[1815]) | ( l_38 [1035] &  i[1815]);
assign l_37[527]    = ( l_38 [1036] & !i[1815]) | ( l_38 [1037] &  i[1815]);
assign l_37[528]    = ( l_38 [1038] & !i[1815]) | ( l_38 [1039] &  i[1815]);
assign l_37[529]    = ( l_38 [1040] & !i[1815]) | ( l_38 [1041] &  i[1815]);
assign l_37[530]    = ( l_38 [1042]);
assign l_37[531]    = ( l_38 [1043]);
assign l_37[532]    = ( l_38 [1044]);
assign l_37[533]    = ( l_38 [1045]);
assign l_37[534]    = ( l_38 [1046]);
assign l_37[535]    = ( l_38 [1047]);
assign l_37[536]    = ( l_38 [1048]);
assign l_37[537]    = ( l_38 [1049]);
assign l_37[538]    = ( l_38 [1050]);
assign l_37[539]    = ( l_38 [1051]);
assign l_37[540]    = ( l_38 [1052]);
assign l_37[541]    = ( l_38 [1053]);
assign l_37[542]    = ( l_38 [1054]);
assign l_37[543]    = ( l_38 [1055]);
assign l_37[544]    = ( l_38 [1056]);
assign l_37[545]    = ( l_38 [1057]);
assign l_37[546]    = ( l_38 [1058]);
assign l_37[547]    = ( l_38 [1059]);
assign l_37[548]    = ( l_38 [1060]);
assign l_37[549]    = ( l_38 [1061]);
assign l_37[550]    = ( l_38 [1062]);
assign l_37[551]    = ( l_38 [1063]);
assign l_37[552]    = ( l_38 [1064]);
assign l_37[553]    = ( l_38 [1065]);
assign l_37[554]    = ( l_38 [1066]);
assign l_37[555]    = ( l_38 [1067]);
assign l_37[556]    = ( l_38 [1068]);
assign l_37[557]    = ( l_38 [1069]);
assign l_37[558]    = ( l_38 [1070]);
assign l_37[559]    = ( l_38 [1071]);
assign l_37[560]    = ( l_38 [1072]);
assign l_37[561]    = ( l_38 [1073]);
assign l_37[562]    = ( l_38 [1074]);
assign l_37[563]    = ( l_38 [1075]);
assign l_37[564]    = ( l_38 [1076]);
assign l_37[565]    = ( l_38 [1077]);
assign l_37[566]    = ( l_38 [1078]);
assign l_37[567]    = ( l_38 [1079]);
assign l_37[568]    = ( l_38 [1080]);
assign l_37[569]    = ( l_38 [1081]);
assign l_37[570]    = ( l_38 [1082]);
assign l_37[571]    = ( l_38 [1083]);
assign l_37[572]    = ( l_38 [1084]);
assign l_37[573]    = ( l_38 [1085]);
assign l_37[574]    = ( l_38 [1086]);
assign l_37[575]    = ( l_38 [1087]);
assign l_37[576]    = ( l_38 [1088]);
assign l_37[577]    = ( l_38 [1089]);
assign l_37[578]    = ( l_38 [1090]);
assign l_37[579]    = ( l_38 [1091]);
assign l_37[580]    = ( l_38 [1092]);
assign l_37[581]    = ( l_38 [1093]);
assign l_37[582]    = ( l_38 [1094]);
assign l_37[583]    = ( l_38 [1095]);
assign l_37[584]    = ( l_38 [1096]);
assign l_37[585]    = ( l_38 [1097]);
assign l_37[586]    = ( l_38 [1098]);
assign l_37[587]    = ( l_38 [1099]);
assign l_37[588]    = ( l_38 [1100]);
assign l_37[589]    = ( l_38 [1101]);
assign l_37[590]    = ( l_38 [1102]);
assign l_37[591]    = ( l_38 [1103]);
assign l_37[592]    = ( l_38 [1104]);
assign l_37[593]    = ( l_38 [1105]);
assign l_37[594]    = ( l_38 [1106]);
assign l_37[595]    = ( l_38 [1107]);
assign l_37[596]    = ( l_38 [1108]);
assign l_37[597]    = ( l_38 [1109]);
assign l_37[598]    = ( l_38 [1110]);
assign l_37[599]    = ( l_38 [1111]);
assign l_37[600]    = ( l_38 [1112]);
assign l_37[601]    = ( l_38 [1113]);
assign l_37[602]    = ( l_38 [1114]);
assign l_37[603]    = ( l_38 [1115]);
assign l_37[604]    = ( l_38 [1116]);
assign l_37[605]    = ( l_38 [1117]);
assign l_37[606]    = ( l_38 [1118]);
assign l_37[607]    = ( l_38 [1119]);
assign l_37[608]    = ( l_38 [1120]);
assign l_37[609]    = ( l_38 [1121]);
assign l_37[610]    = ( l_38 [1122]);
assign l_37[611]    = ( l_38 [1123]);
assign l_37[612]    = ( l_38 [1124]);
assign l_37[613]    = ( l_38 [1125]);
assign l_37[614]    = ( l_38 [1126]);
assign l_37[615]    = ( l_38 [1127]);
assign l_37[616]    = ( l_38 [1128]);
assign l_37[617]    = ( l_38 [1129]);
assign l_37[618]    = ( l_38 [1130]);
assign l_37[619]    = ( l_38 [1131]);
assign l_37[620]    = ( l_38 [1132]);
assign l_37[621]    = ( l_38 [1133]);
assign l_37[622]    = ( l_38 [1134]);
assign l_37[623]    = ( l_38 [1135]);
assign l_37[624]    = ( l_38 [1136]);
assign l_37[625]    = ( l_38 [1137]);
assign l_37[626]    = ( l_38 [1138]);
assign l_37[627]    = ( l_38 [1139]);
assign l_37[628]    = ( l_38 [1140]);
assign l_37[629]    = ( l_38 [1141]);
assign l_37[630]    = ( l_38 [1142]);
assign l_37[631]    = ( l_38 [1143]);
assign l_37[632]    = ( l_38 [1144]);
assign l_37[633]    = ( l_38 [1145]);
assign l_37[634]    = ( l_38 [1146]);
assign l_37[635]    = ( l_38 [1147]);
assign l_37[636]    = ( l_38 [1148]);
assign l_37[637]    = ( l_38 [1149]);
assign l_37[638]    = ( l_38 [1150]);
assign l_37[639]    = ( l_38 [1151]);
assign l_37[640]    = ( l_38 [1152]);
assign l_37[641]    = ( l_38 [1153]);
assign l_37[642]    = ( l_38 [1154]);
assign l_37[643]    = ( l_38 [1155]);
assign l_37[644]    = ( l_38 [1156]);
assign l_37[645]    = ( l_38 [1157]);
assign l_37[646]    = ( l_38 [1158]);
assign l_37[647]    = ( l_38 [1159]);
assign l_37[648]    = ( l_38 [1160]);
assign l_37[649]    = ( l_38 [1161]);
assign l_37[650]    = ( l_38 [1162]);
assign l_37[651]    = ( l_38 [1163]);
assign l_37[652]    = ( l_38 [1164]);
assign l_37[653]    = ( l_38 [1165]);
assign l_37[654]    = ( l_38 [1166]);
assign l_37[655]    = ( l_38 [1167]);
assign l_37[656]    = ( l_38 [1168]);
assign l_37[657]    = ( l_38 [1169]);
assign l_37[658]    = ( l_38 [1170]);
assign l_37[659]    = ( l_38 [1171]);
assign l_37[660]    = ( l_38 [1172]);
assign l_37[661]    = ( l_38 [1173]);
assign l_37[662]    = ( l_38 [1174]);
assign l_37[663]    = ( l_38 [1175]);
assign l_37[664]    = ( l_38 [1176]);
assign l_37[665]    = ( l_38 [1177]);
assign l_37[666]    = ( l_38 [1178]);
assign l_37[667]    = ( l_38 [1179]);
assign l_37[668]    = ( l_38 [1180]);
assign l_37[669]    = ( l_38 [1181]);
assign l_37[670]    = ( l_38 [1182]);
assign l_37[671]    = ( l_38 [1183]);
assign l_37[672]    = ( l_38 [1184]);
assign l_37[673]    = ( l_38 [1185]);
assign l_37[674]    = ( l_38 [1186]);
assign l_37[675]    = ( l_38 [1187]);
assign l_37[676]    = ( l_38 [1188]);
assign l_37[677]    = ( l_38 [1189]);
assign l_37[678]    = ( l_38 [1190]);
assign l_37[679]    = ( l_38 [1191]);
assign l_37[680]    = ( l_38 [1192]);
assign l_37[681]    = ( l_38 [1193]);
assign l_37[682]    = ( l_38 [1194]);
assign l_37[683]    = ( l_38 [1195]);
assign l_37[684]    = ( l_38 [1196]);
assign l_37[685]    = ( l_38 [1197]);
assign l_37[686]    = ( l_38 [1198]);
assign l_37[687]    = ( l_38 [1199]);
assign l_37[688]    = ( l_38 [1200]);
assign l_37[689]    = ( l_38 [1201]);
assign l_37[690]    = ( l_38 [1202]);
assign l_37[691]    = ( l_38 [1203]);
assign l_37[692]    = ( l_38 [1204]);
assign l_37[693]    = ( l_38 [1205]);
assign l_37[694]    = ( l_38 [1206]);
assign l_37[695]    = ( l_38 [1207]);
assign l_37[696]    = ( l_38 [1208]);
assign l_37[697]    = ( l_38 [1209]);
assign l_37[698]    = ( l_38 [1210]);
assign l_37[699]    = ( l_38 [1211]);
assign l_37[700]    = ( l_38 [1212]);
assign l_37[701]    = ( l_38 [1213]);
assign l_37[702]    = ( l_38 [1214]);
assign l_37[703]    = ( l_38 [1215]);
assign l_37[704]    = ( l_38 [1216]);
assign l_37[705]    = ( l_38 [1217]);
assign l_37[706]    = ( l_38 [1218]);
assign l_37[707]    = ( l_38 [1219]);
assign l_37[708]    = ( l_38 [1220]);
assign l_37[709]    = ( l_38 [1221]);
assign l_37[710]    = ( l_38 [1222]);
assign l_37[711]    = ( l_38 [1223]);
assign l_37[712]    = ( l_38 [1224]);
assign l_37[713]    = ( l_38 [1225]);
assign l_37[714]    = ( l_38 [1226]);
assign l_37[715]    = ( l_38 [1227]);
assign l_37[716]    = ( l_38 [1228]);
assign l_37[717]    = ( l_38 [1229]);
assign l_37[718]    = ( l_38 [1230]);
assign l_37[719]    = ( l_38 [1231]);
assign l_37[720]    = ( l_38 [1232]);
assign l_37[721]    = ( l_38 [1233]);
assign l_37[722]    = ( l_38 [1234]);
assign l_37[723]    = ( l_38 [1235]);
assign l_37[724]    = ( l_38 [1236]);
assign l_37[725]    = ( l_38 [1237]);
assign l_37[726]    = ( l_38 [1238]);
assign l_37[727]    = ( l_38 [1239]);
assign l_37[728]    = ( l_38 [1240]);
assign l_37[729]    = ( l_38 [1241]);
assign l_37[730]    = ( l_38 [1242]);
assign l_37[731]    = ( l_38 [1243]);
assign l_37[732]    = ( l_38 [1244]);
assign l_37[733]    = ( l_38 [1245]);
assign l_37[734]    = ( l_38 [1246]);
assign l_37[735]    = ( l_38 [1247]);
assign l_37[736]    = ( l_38 [1248]);
assign l_37[737]    = ( l_38 [1249]);
assign l_37[738]    = ( l_38 [1250]);
assign l_37[739]    = ( l_38 [1251]);
assign l_37[740]    = ( l_38 [1252]);
assign l_37[741]    = ( l_38 [1253]);
assign l_37[742]    = ( l_38 [1254]);
assign l_37[743]    = ( l_38 [1255]);
assign l_37[744]    = ( l_38 [1256]);
assign l_37[745]    = ( l_38 [1257]);
assign l_37[746]    = ( l_38 [1258]);
assign l_37[747]    = ( l_38 [1259]);
assign l_37[748]    = ( l_38 [1260]);
assign l_37[749]    = ( l_38 [1261]);
assign l_37[750]    = ( l_38 [1262]);
assign l_37[751]    = ( l_38 [1263]);
assign l_37[752]    = ( l_38 [1264]);
assign l_37[753]    = ( l_38 [1265]);
assign l_37[754]    = ( l_38 [1266]);
assign l_37[755]    = ( l_38 [1267]);
assign l_37[756]    = ( l_38 [1268]);
assign l_37[757]    = ( l_38 [1269]);
assign l_37[758]    = ( l_38 [1270]);
assign l_37[759]    = ( l_38 [1271]);
assign l_37[760]    = ( l_38 [1272]);
assign l_37[761]    = ( l_38 [1273]);
assign l_37[762]    = ( l_38 [1274]);
assign l_37[763]    = ( l_38 [1275]);
assign l_37[764]    = ( l_38 [1276]);
assign l_37[765]    = ( l_38 [1277]);
assign l_37[766]    = ( l_38 [1278]);
assign l_37[767]    = ( l_38 [1279]);
assign l_37[768]    = ( l_38 [1280]);
assign l_37[769]    = ( l_38 [1281]);
assign l_37[770]    = ( l_38 [1282]);
assign l_37[771]    = ( l_38 [1283]);
assign l_37[772]    = ( l_38 [1284]);
assign l_37[773]    = ( l_38 [1285]);
assign l_37[774]    = ( l_38 [1286]);
assign l_37[775]    = ( l_38 [1287]);
assign l_37[776]    = ( l_38 [1288]);
assign l_37[777]    = ( l_38 [1289]);
assign l_37[778]    = ( l_38 [1290]);
assign l_37[779]    = ( l_38 [1291]);
assign l_37[780]    = ( l_38 [1292]);
assign l_37[781]    = ( l_38 [1293]);
assign l_37[782]    = ( l_38 [1294]);
assign l_37[783]    = ( l_38 [1295]);
assign l_37[784]    = ( l_38 [1296]);
assign l_37[785]    = ( l_38 [1297]);
assign l_37[786]    = ( l_38 [1298]);
assign l_37[787]    = ( l_38 [1299]);
assign l_37[788]    = ( l_38 [1300]);
assign l_37[789]    = ( l_38 [1301]);
assign l_37[790]    = ( l_38 [1302]);
assign l_37[791]    = ( l_38 [1303]);
assign l_37[792]    = ( l_38 [1304]);
assign l_37[793]    = ( l_38 [1305]);
assign l_37[794]    = ( l_38 [1306]);
assign l_37[795]    = ( l_38 [1307]);
assign l_37[796]    = ( l_38 [1308]);
assign l_37[797]    = ( l_38 [1309]);
assign l_37[798]    = ( l_38 [1310]);
assign l_37[799]    = ( l_38 [1311]);
assign l_37[800]    = ( l_38 [1312]);
assign l_37[801]    = ( l_38 [1313]);
assign l_37[802]    = ( l_38 [1314]);
assign l_37[803]    = ( l_38 [1315]);
assign l_37[804]    = ( l_38 [1316]);
assign l_37[805]    = ( l_38 [1317]);
assign l_37[806]    = ( l_38 [1318]);
assign l_37[807]    = ( l_38 [1319]);
assign l_37[808]    = ( l_38 [1320]);
assign l_37[809]    = ( l_38 [1321]);
assign l_37[810]    = ( l_38 [1322]);
assign l_37[811]    = ( l_38 [1323]);
assign l_37[812]    = ( l_38 [1324]);
assign l_37[813]    = ( l_38 [1325]);
assign l_37[814]    = ( l_38 [1326]);
assign l_37[815]    = ( l_38 [1327]);
assign l_37[816]    = ( l_38 [1328]);
assign l_37[817]    = ( l_38 [1329]);
assign l_37[818]    = ( l_38 [1330]);
assign l_37[819]    = ( l_38 [1331]);
assign l_37[820]    = ( l_38 [1332]);
assign l_37[821]    = ( l_38 [1333]);
assign l_37[822]    = ( l_38 [1334]);
assign l_37[823]    = ( l_38 [1335]);
assign l_37[824]    = ( l_38 [1336]);
assign l_37[825]    = ( l_38 [1337]);
assign l_37[826]    = ( l_38 [1338]);
assign l_37[827]    = ( l_38 [1339]);
assign l_37[828]    = ( l_38 [1340]);
assign l_37[829]    = ( l_38 [1341]);
assign l_37[830]    = ( l_38 [1342]);
assign l_37[831]    = ( l_38 [1343]);
assign l_37[832]    = ( l_38 [1344]);
assign l_37[833]    = ( l_38 [1345]);
assign l_37[834]    = ( l_38 [1346]);
assign l_37[835]    = ( l_38 [1347]);
assign l_37[836]    = ( l_38 [1348]);
assign l_37[837]    = ( l_38 [1349]);
assign l_37[838]    = ( l_38 [1350]);
assign l_37[839]    = ( l_38 [1351]);
assign l_37[840]    = ( l_38 [1352]);
assign l_37[841]    = ( l_38 [1353]);
assign l_37[842]    = ( l_38 [1354]);
assign l_37[843]    = ( l_38 [1355]);
assign l_37[844]    = ( l_38 [1356]);
assign l_37[845]    = ( l_38 [1357]);
assign l_37[846]    = ( l_38 [1358]);
assign l_37[847]    = ( l_38 [1359]);
assign l_37[848]    = ( l_38 [1360]);
assign l_37[849]    = ( l_38 [1361]);
assign l_37[850]    = ( l_38 [1362]);
assign l_37[851]    = ( l_38 [1363]);
assign l_37[852]    = ( l_38 [1364]);
assign l_37[853]    = ( l_38 [1365]);
assign l_37[854]    = ( l_38 [1366]);
assign l_37[855]    = ( l_38 [1367]);
assign l_37[856]    = ( l_38 [1368]);
assign l_37[857]    = ( l_38 [1369]);
assign l_37[858]    = ( l_38 [1370]);
assign l_37[859]    = ( l_38 [1371]);
assign l_37[860]    = ( l_38 [1372]);
assign l_37[861]    = ( l_38 [1373]);
assign l_37[862]    = ( l_38 [1374]);
assign l_37[863]    = ( l_38 [1375]);
assign l_37[864]    = ( l_38 [1376]);
assign l_37[865]    = ( l_38 [1377]);
assign l_37[866]    = ( l_38 [1378]);
assign l_37[867]    = ( l_38 [1379]);
assign l_37[868]    = ( l_38 [1380]);
assign l_37[869]    = ( l_38 [1381]);
assign l_37[870]    = ( l_38 [1382]);
assign l_37[871]    = ( l_38 [1383]);
assign l_37[872]    = ( l_38 [1384]);
assign l_37[873]    = ( l_38 [1385]);
assign l_37[874]    = ( l_38 [1386]);
assign l_37[875]    = ( l_38 [1387]);
assign l_37[876]    = ( l_38 [1388]);
assign l_37[877]    = ( l_38 [1389]);
assign l_37[878]    = ( l_38 [1390]);
assign l_37[879]    = ( l_38 [1391]);
assign l_37[880]    = ( l_38 [1392]);
assign l_37[881]    = ( l_38 [1393]);
assign l_37[882]    = ( l_38 [1394]);
assign l_37[883]    = ( l_38 [1395]);
assign l_37[884]    = ( l_38 [1396]);
assign l_37[885]    = ( l_38 [1397]);
assign l_37[886]    = ( l_38 [1398]);
assign l_37[887]    = ( l_38 [1399]);
assign l_37[888]    = ( l_38 [1400]);
assign l_37[889]    = ( l_38 [1401]);
assign l_37[890]    = ( l_38 [1402]);
assign l_37[891]    = ( l_38 [1403]);
assign l_37[892]    = ( l_38 [1404]);
assign l_37[893]    = ( l_38 [1405]);
assign l_37[894]    = ( l_38 [1406]);
assign l_37[895]    = ( l_38 [1407]);
assign l_37[896]    = ( l_38 [1408]);
assign l_37[897]    = ( l_38 [1409]);
assign l_37[898]    = ( l_38 [1410]);
assign l_37[899]    = ( l_38 [1411]);
assign l_37[900]    = ( l_38 [1412]);
assign l_37[901]    = ( l_38 [1413]);
assign l_37[902]    = ( l_38 [1414]);
assign l_37[903]    = ( l_38 [1415]);
assign l_37[904]    = ( l_38 [1416]);
assign l_37[905]    = ( l_38 [1417]);
assign l_37[906]    = ( l_38 [1418]);
assign l_37[907]    = ( l_38 [1419]);
assign l_37[908]    = ( l_38 [1420]);
assign l_37[909]    = ( l_38 [1421]);
assign l_37[910]    = ( l_38 [1422]);
assign l_37[911]    = ( l_38 [1423]);
assign l_37[912]    = ( l_38 [1424]);
assign l_37[913]    = ( l_38 [1425]);
assign l_37[914]    = ( l_38 [1426]);
assign l_37[915]    = ( l_38 [1427]);
assign l_37[916]    = ( l_38 [1428]);
assign l_37[917]    = ( l_38 [1429]);
assign l_37[918]    = ( l_38 [1430]);
assign l_37[919]    = ( l_38 [1431]);
assign l_37[920]    = ( l_38 [1432]);
assign l_37[921]    = ( l_38 [1433]);
assign l_37[922]    = ( l_38 [1434]);
assign l_37[923]    = ( l_38 [1435]);
assign l_37[924]    = ( l_38 [1436]);
assign l_37[925]    = ( l_38 [1437]);
assign l_37[926]    = ( l_38 [1438]);
assign l_37[927]    = ( l_38 [1439]);
assign l_37[928]    = ( l_38 [1440]);
assign l_37[929]    = ( l_38 [1441]);
assign l_37[930]    = ( l_38 [1442]);
assign l_37[931]    = ( l_38 [1443]);
assign l_37[932]    = ( l_38 [1444]);
assign l_37[933]    = ( l_38 [1445]);
assign l_37[934]    = ( l_38 [1446]);
assign l_37[935]    = ( l_38 [1447]);
assign l_37[936]    = ( l_38 [1448]);
assign l_37[937]    = ( l_38 [1449]);
assign l_37[938]    = ( l_38 [1450]);
assign l_37[939]    = ( l_38 [1451]);
assign l_37[940]    = ( l_38 [1452]);
assign l_37[941]    = ( l_38 [1453]);
assign l_37[942]    = ( l_38 [1454]);
assign l_37[943]    = ( l_38 [1455]);
assign l_37[944]    = ( l_38 [1456]);
assign l_37[945]    = ( l_38 [1457]);
assign l_37[946]    = ( l_38 [1458]);
assign l_37[947]    = ( l_38 [1459]);
assign l_37[948]    = ( l_38 [1460]);
assign l_37[949]    = ( l_38 [1461]);
assign l_37[950]    = ( l_38 [1462]);
assign l_37[951]    = ( l_38 [1463]);
assign l_37[952]    = ( l_38 [1464]);
assign l_37[953]    = ( l_38 [1465]);
assign l_37[954]    = ( l_38 [1466]);
assign l_37[955]    = ( l_38 [1467]);
assign l_37[956]    = ( l_38 [1468]);
assign l_37[957]    = ( l_38 [1469]);
assign l_37[958]    = ( l_38 [1470]);
assign l_37[959]    = ( l_38 [1471]);
assign l_37[960]    = ( l_38 [1472]);
assign l_37[961]    = ( l_38 [1473]);
assign l_37[962]    = ( l_38 [1474]);
assign l_37[963]    = ( l_38 [1475]);
assign l_37[964]    = ( l_38 [1476]);
assign l_37[965]    = ( l_38 [1477]);
assign l_37[966]    = ( l_38 [1478]);
assign l_37[967]    = ( l_38 [1479]);
assign l_37[968]    = ( l_38 [1480]);
assign l_37[969]    = ( l_38 [1481]);
assign l_37[970]    = ( l_38 [1482]);
assign l_37[971]    = ( l_38 [1483]);
assign l_37[972]    = ( l_38 [1484]);
assign l_37[973]    = ( l_38 [1485]);
assign l_37[974]    = ( l_38 [1486]);
assign l_37[975]    = ( l_38 [1487]);
assign l_37[976]    = ( l_38 [1488]);
assign l_37[977]    = ( l_38 [1489]);
assign l_37[978]    = ( l_38 [1490]);
assign l_37[979]    = ( l_38 [1491]);
assign l_37[980]    = ( l_38 [1492]);
assign l_37[981]    = ( l_38 [1493]);
assign l_37[982]    = ( l_38 [1494]);
assign l_37[983]    = ( l_38 [1495]);
assign l_37[984]    = ( l_38 [1496]);
assign l_37[985]    = ( l_38 [1497]);
assign l_37[986]    = ( l_38 [1498]);
assign l_37[987]    = ( l_38 [1499]);
assign l_37[988]    = ( l_38 [1500]);
assign l_37[989]    = ( l_38 [1501]);
assign l_37[990]    = ( l_38 [1502]);
assign l_37[991]    = ( l_38 [1503]);
assign l_37[992]    = ( l_38 [1504]);
assign l_37[993]    = ( l_38 [1505]);
assign l_37[994]    = ( l_38 [1506]);
assign l_37[995]    = ( l_38 [1507]);
assign l_37[996]    = ( l_38 [1508]);
assign l_37[997]    = ( l_38 [1509]);
assign l_37[998]    = ( l_38 [1510]);
assign l_37[999]    = ( l_38 [1511]);
assign l_37[1000]    = ( l_38 [1512]);
assign l_37[1001]    = ( l_38 [1513]);
assign l_37[1002]    = ( l_38 [1514]);
assign l_37[1003]    = ( l_38 [1515]);
assign l_37[1004]    = ( l_38 [1516]);
assign l_37[1005]    = ( l_38 [1517]);
assign l_37[1006]    = ( l_38 [1518]);
assign l_37[1007]    = ( l_38 [1519]);
assign l_37[1008]    = ( l_38 [1520]);
assign l_37[1009]    = ( l_38 [1521]);
assign l_37[1010]    = ( l_38 [1522]);
assign l_37[1011]    = ( l_38 [1523]);
assign l_37[1012]    = ( l_38 [1524]);
assign l_37[1013]    = ( l_38 [1525]);
assign l_37[1014]    = ( l_38 [1526]);
assign l_37[1015]    = ( l_38 [1527]);
assign l_37[1016]    = ( l_38 [1528]);
assign l_37[1017]    = ( l_38 [1529]);
assign l_37[1018]    = ( l_38 [1530]);
assign l_37[1019]    = ( l_38 [1531]);
assign l_37[1020]    = ( l_38 [1532]);
assign l_37[1021]    = ( l_38 [1533]);
assign l_37[1022]    = ( l_38 [1534]);
assign l_37[1023]    = ( l_38 [1535]);
assign l_37[1024]    = ( l_38 [1536]);
assign l_37[1025]    = ( l_38 [1537]);
assign l_37[1026]    = ( l_38 [1538]);
assign l_37[1027]    = ( l_38 [1539]);
assign l_37[1028]    = ( l_38 [1540]);
assign l_37[1029]    = ( l_38 [1541]);
assign l_37[1030]    = ( l_38 [1542]);
assign l_37[1031]    = ( l_38 [1543]);
assign l_37[1032]    = ( l_38 [1544]);
assign l_37[1033]    = ( l_38 [1545]);
assign l_37[1034]    = ( l_38 [1546]);
assign l_37[1035]    = ( l_38 [1547]);
assign l_37[1036]    = ( l_38 [1548]);
assign l_37[1037]    = ( l_38 [1549]);
assign l_37[1038]    = ( l_38 [1550]);
assign l_37[1039]    = ( l_38 [1551]);
assign l_37[1040]    = ( l_38 [1552]);
assign l_37[1041]    = ( l_38 [1553]);
assign l_37[1042]    = ( l_38 [1554]);
assign l_37[1043]    = ( l_38 [1555]);
assign l_37[1044]    = ( l_38 [1556]);
assign l_37[1045]    = ( l_38 [1557]);
assign l_37[1046]    = ( l_38 [1558]);
assign l_37[1047]    = ( l_38 [1559]);
assign l_37[1048]    = ( l_38 [1560]);
assign l_37[1049]    = ( l_38 [1561]);
assign l_37[1050]    = ( l_38 [1562]);
assign l_37[1051]    = ( l_38 [1563]);
assign l_37[1052]    = ( l_38 [1564]);
assign l_37[1053]    = ( l_38 [1565]);
assign l_37[1054]    = ( l_38 [1566]);
assign l_37[1055]    = ( l_38 [1567]);
assign l_37[1056]    = ( l_38 [1568]);
assign l_37[1057]    = ( l_38 [1569]);
assign l_37[1058]    = ( l_38 [1570]);
assign l_37[1059]    = ( l_38 [1571]);
assign l_37[1060]    = ( l_38 [1572]);
assign l_37[1061]    = ( l_38 [1573]);
assign l_37[1062]    = ( l_38 [1574]);
assign l_37[1063]    = ( l_38 [1575]);
assign l_37[1064]    = ( l_38 [1576]);
assign l_37[1065]    = ( l_38 [1577]);
assign l_37[1066]    = ( l_38 [1578]);
assign l_37[1067]    = ( l_38 [1579]);
assign l_37[1068]    = ( l_38 [1580]);
assign l_37[1069]    = ( l_38 [1581]);
assign l_37[1070]    = ( l_38 [1582]);
assign l_37[1071]    = ( l_38 [1583]);
assign l_37[1072]    = ( l_38 [1584]);
assign l_37[1073]    = ( l_38 [1585]);
assign l_37[1074]    = ( l_38 [1586]);
assign l_37[1075]    = ( l_38 [1587]);
assign l_37[1076]    = ( l_38 [1588]);
assign l_37[1077]    = ( l_38 [1589]);
assign l_37[1078]    = ( l_38 [1590]);
assign l_37[1079]    = ( l_38 [1591]);
assign l_37[1080]    = ( l_38 [1592]);
assign l_37[1081]    = ( l_38 [1593]);
assign l_37[1082]    = ( l_38 [1594]);
assign l_37[1083]    = ( l_38 [1595]);
assign l_37[1084]    = ( l_38 [1596]);
assign l_37[1085]    = ( l_38 [1597]);
assign l_37[1086]    = ( l_38 [1598]);
assign l_37[1087]    = ( l_38 [1599]);
assign l_37[1088]    = ( l_38 [1600]);
assign l_37[1089]    = ( l_38 [1601]);
assign l_37[1090]    = ( l_38 [1602]);
assign l_37[1091]    = ( l_38 [1603]);
assign l_37[1092]    = ( l_38 [1604]);
assign l_37[1093]    = ( l_38 [1605]);
assign l_37[1094]    = ( l_38 [1606]);
assign l_37[1095]    = ( l_38 [1607]);
assign l_37[1096]    = ( l_38 [1608]);
assign l_37[1097]    = ( l_38 [1609]);
assign l_37[1098]    = ( l_38 [1610]);
assign l_37[1099]    = ( l_38 [1611]);
assign l_37[1100]    = ( l_38 [1612]);
assign l_37[1101]    = ( l_38 [1613]);
assign l_37[1102]    = ( l_38 [1614]);
assign l_37[1103]    = ( l_38 [1615]);
assign l_37[1104]    = ( l_38 [1616]);
assign l_37[1105]    = ( l_38 [1617]);
assign l_37[1106]    = ( l_38 [1618]);
assign l_37[1107]    = ( l_38 [1619]);
assign l_37[1108]    = ( l_38 [1620]);
assign l_37[1109]    = ( l_38 [1621]);
assign l_37[1110]    = ( l_38 [1622]);
assign l_37[1111]    = ( l_38 [1623]);
assign l_37[1112]    = ( l_38 [1624]);
assign l_37[1113]    = ( l_38 [1625]);
assign l_37[1114]    = ( l_38 [1626]);
assign l_37[1115]    = ( l_38 [1627]);
assign l_37[1116]    = ( l_38 [1628]);
assign l_37[1117]    = ( l_38 [1629]);
assign l_37[1118]    = ( l_38 [1630]);
assign l_37[1119]    = ( l_38 [1631]);
assign l_37[1120]    = ( l_38 [1632]);
assign l_37[1121]    = ( l_38 [1633]);
assign l_37[1122]    = ( l_38 [1634]);
assign l_37[1123]    = ( l_38 [1635]);
assign l_37[1124]    = ( l_38 [1636]);
assign l_37[1125]    = ( l_38 [1637]);
assign l_37[1126]    = ( l_38 [1638]);
assign l_37[1127]    = ( l_38 [1639]);
assign l_37[1128]    = ( l_38 [1640]);
assign l_37[1129]    = ( l_38 [1641]);
assign l_37[1130]    = ( l_38 [1642]);
assign l_37[1131]    = ( l_38 [1643]);
assign l_37[1132]    = ( l_38 [1644]);
assign l_37[1133]    = ( l_38 [1645]);
assign l_37[1134]    = ( l_38 [1646]);
assign l_37[1135]    = ( l_38 [1647]);
assign l_37[1136]    = ( l_38 [1648]);
assign l_37[1137]    = ( l_38 [1649]);
assign l_37[1138]    = ( l_38 [1650]);
assign l_37[1139]    = ( l_38 [1651]);
assign l_37[1140]    = ( l_38 [1652]);
assign l_37[1141]    = ( l_38 [1653]);
assign l_37[1142]    = ( l_38 [1654]);
assign l_37[1143]    = ( l_38 [1655]);
assign l_37[1144]    = ( l_38 [1656]);
assign l_37[1145]    = ( l_38 [1657]);
assign l_37[1146]    = ( l_38 [1658]);
assign l_37[1147]    = ( l_38 [1659]);
assign l_37[1148]    = ( l_38 [1660]);
assign l_37[1149]    = ( l_38 [1661]);
assign l_37[1150]    = ( l_38 [1662]);
assign l_37[1151]    = ( l_38 [1663]);
assign l_37[1152]    = ( l_38 [1664]);
assign l_37[1153]    = ( l_38 [1665]);
assign l_37[1154]    = ( l_38 [1666]);
assign l_37[1155]    = ( l_38 [1667]);
assign l_37[1156]    = ( l_38 [1668]);
assign l_37[1157]    = ( l_38 [1669]);
assign l_37[1158]    = ( l_38 [1670]);
assign l_37[1159]    = ( l_38 [1671]);
assign l_37[1160]    = ( l_38 [1672]);
assign l_37[1161]    = ( l_38 [1673]);
assign l_37[1162]    = ( l_38 [1674]);
assign l_37[1163]    = ( l_38 [1675]);
assign l_37[1164]    = ( l_38 [1676]);
assign l_37[1165]    = ( l_38 [1677]);
assign l_37[1166]    = ( l_38 [1678]);
assign l_37[1167]    = ( l_38 [1679]);
assign l_37[1168]    = ( l_38 [1680]);
assign l_37[1169]    = ( l_38 [1681]);
assign l_37[1170]    = ( l_38 [1682]);
assign l_37[1171]    = ( l_38 [1683]);
assign l_37[1172]    = ( l_38 [1684]);
assign l_37[1173]    = ( l_38 [1685]);
assign l_37[1174]    = ( l_38 [1686]);
assign l_37[1175]    = ( l_38 [1687]);
assign l_37[1176]    = ( l_38 [1688]);
assign l_37[1177]    = ( l_38 [1689]);
assign l_37[1178]    = ( l_38 [1690]);
assign l_37[1179]    = ( l_38 [1691]);
assign l_37[1180]    = ( l_38 [1692]);
assign l_37[1181]    = ( l_38 [1693]);
assign l_37[1182]    = ( l_38 [1694]);
assign l_37[1183]    = ( l_38 [1695]);
assign l_37[1184]    = ( l_38 [1696]);
assign l_37[1185]    = ( l_38 [1697]);
assign l_37[1186]    = ( l_38 [1698]);
assign l_37[1187]    = ( l_38 [1699]);
assign l_37[1188]    = ( l_38 [1700]);
assign l_37[1189]    = ( l_38 [1701]);
assign l_37[1190]    = ( l_38 [1702]);
assign l_37[1191]    = ( l_38 [1703]);
assign l_37[1192]    = ( l_38 [1704]);
assign l_37[1193]    = ( l_38 [1705]);
assign l_37[1194]    = ( l_38 [1706]);
assign l_37[1195]    = ( l_38 [1707]);
assign l_37[1196]    = ( l_38 [1708]);
assign l_37[1197]    = ( l_38 [1709]);
assign l_37[1198]    = ( l_38 [1710]);
assign l_37[1199]    = ( l_38 [1711]);
assign l_37[1200]    = ( l_38 [1712]);
assign l_37[1201]    = ( l_38 [1713]);
assign l_37[1202]    = ( l_38 [1714]);
assign l_37[1203]    = ( l_38 [1715]);
assign l_37[1204]    = ( l_38 [1716]);
assign l_37[1205]    = ( l_38 [1717]);
assign l_37[1206]    = ( l_38 [1718]);
assign l_37[1207]    = ( l_38 [1719]);
assign l_37[1208]    = ( l_38 [1720]);
assign l_37[1209]    = ( l_38 [1721]);
assign l_37[1210]    = ( l_38 [1722]);
assign l_37[1211]    = ( l_38 [1723]);
assign l_37[1212]    = ( l_38 [1724]);
assign l_37[1213]    = ( l_38 [1725]);
assign l_37[1214]    = ( l_38 [1726]);
assign l_37[1215]    = ( l_38 [1727]);
assign l_37[1216]    = ( l_38 [1728]);
assign l_37[1217]    = ( l_38 [1729]);
assign l_37[1218]    = ( l_38 [1730]);
assign l_37[1219]    = ( l_38 [1731]);
assign l_37[1220]    = ( l_38 [1732]);
assign l_37[1221]    = ( l_38 [1733]);
assign l_37[1222]    = ( l_38 [1734]);
assign l_37[1223]    = ( l_38 [1735]);
assign l_37[1224]    = ( l_38 [1736]);
assign l_37[1225]    = ( l_38 [1737]);
assign l_37[1226]    = ( l_38 [1738]);
assign l_37[1227]    = ( l_38 [1739]);
assign l_37[1228]    = ( l_38 [1740]);
assign l_37[1229]    = ( l_38 [1741]);
assign l_37[1230]    = ( l_38 [1742]);
assign l_37[1231]    = ( l_38 [1743]);
assign l_37[1232]    = ( l_38 [1744]);
assign l_37[1233]    = ( l_38 [1745]);
assign l_37[1234]    = ( l_38 [1746]);
assign l_37[1235]    = ( l_38 [1747]);
assign l_37[1236]    = ( l_38 [1748]);
assign l_37[1237]    = ( l_38 [1749]);
assign l_37[1238]    = ( l_38 [1750]);
assign l_37[1239]    = ( l_38 [1751]);
assign l_37[1240]    = ( l_38 [1752]);
assign l_37[1241]    = ( l_38 [1753]);
assign l_37[1242]    = ( l_38 [1754]);
assign l_37[1243]    = ( l_38 [1755]);
assign l_37[1244]    = ( l_38 [1756]);
assign l_37[1245]    = ( l_38 [1757]);
assign l_37[1246]    = ( l_38 [1758]);
assign l_37[1247]    = ( l_38 [1759]);
assign l_37[1248]    = ( l_38 [1760]);
assign l_37[1249]    = ( l_38 [1761]);
assign l_37[1250]    = ( l_38 [1762]);
assign l_37[1251]    = ( l_38 [1763]);
assign l_37[1252]    = ( l_38 [1764]);
assign l_37[1253]    = ( l_38 [1765]);
assign l_37[1254]    = ( l_38 [1766]);
assign l_37[1255]    = ( l_38 [1767]);
assign l_37[1256]    = ( l_38 [1768]);
assign l_37[1257]    = ( l_38 [1769]);
assign l_37[1258]    = ( l_38 [1770]);
assign l_37[1259]    = ( l_38 [1771]);
assign l_37[1260]    = ( l_38 [1772]);
assign l_37[1261]    = ( l_38 [1773]);
assign l_37[1262]    = ( l_38 [1774]);
assign l_37[1263]    = ( l_38 [1775]);
assign l_37[1264]    = ( l_38 [1776]);
assign l_37[1265]    = ( l_38 [1777]);
assign l_37[1266]    = ( l_38 [1778]);
assign l_37[1267]    = ( l_38 [1779]);
assign l_37[1268]    = ( l_38 [1780]);
assign l_37[1269]    = ( l_38 [1781]);
assign l_37[1270]    = ( l_38 [1782]);
assign l_37[1271]    = ( l_38 [1783]);
assign l_37[1272]    = ( l_38 [1784]);
assign l_37[1273]    = ( l_38 [1785]);
assign l_37[1274]    = ( l_38 [1786]);
assign l_37[1275]    = ( l_38 [1787]);
assign l_37[1276]    = ( l_38 [1788]);
assign l_37[1277]    = ( l_38 [1789]);
assign l_37[1278]    = ( l_38 [1790]);
assign l_37[1279]    = ( l_38 [1791]);
assign l_37[1280]    = ( l_38 [1792]);
assign l_37[1281]    = ( l_38 [1793]);
assign l_37[1282]    = ( l_38 [1794]);
assign l_37[1283]    = ( l_38 [1795]);
assign l_37[1284]    = ( l_38 [1796]);
assign l_37[1285]    = ( l_38 [1797]);
assign l_37[1286]    = ( l_38 [1798]);
assign l_37[1287]    = ( l_38 [1799]);
assign l_37[1288]    = ( l_38 [1800]);
assign l_37[1289]    = ( l_38 [1801]);
assign l_37[1290]    = ( l_38 [1802]);
assign l_37[1291]    = ( l_38 [1803]);
assign l_37[1292]    = ( l_38 [1804]);
assign l_37[1293]    = ( l_38 [1805]);
assign l_37[1294]    = ( l_38 [1806]);
assign l_37[1295]    = ( l_38 [1807]);
assign l_37[1296]    = ( l_38 [1808]);
assign l_37[1297]    = ( l_38 [1809]);
assign l_37[1298]    = ( l_38 [1810]);
assign l_37[1299]    = ( l_38 [1811]);
assign l_37[1300]    = ( l_38 [1812]);
assign l_37[1301]    = ( l_38 [1813]);
assign l_37[1302]    = ( l_38 [1814]);
assign l_37[1303]    = ( l_38 [1815]);
assign l_37[1304]    = ( l_38 [1816]);
assign l_37[1305]    = ( l_38 [1817]);
assign l_37[1306]    = ( l_38 [1818]);
assign l_37[1307]    = ( l_38 [1819]);
assign l_37[1308]    = ( l_38 [1820]);
assign l_37[1309]    = ( l_38 [1821]);
assign l_37[1310]    = ( l_38 [1822]);
assign l_37[1311]    = ( l_38 [1823]);
assign l_37[1312]    = ( l_38 [1824]);
assign l_37[1313]    = ( l_38 [1825]);
assign l_37[1314]    = ( l_38 [1826]);
assign l_37[1315]    = ( l_38 [1827]);
assign l_37[1316]    = ( l_38 [1828]);
assign l_37[1317]    = ( l_38 [1829]);
assign l_37[1318]    = ( l_38 [1830]);
assign l_37[1319]    = ( l_38 [1831]);
assign l_37[1320]    = ( l_38 [1832]);
assign l_37[1321]    = ( l_38 [1833]);
assign l_37[1322]    = ( l_38 [1834]);
assign l_37[1323]    = ( l_38 [1835]);
assign l_37[1324]    = ( l_38 [1836]);
assign l_37[1325]    = ( l_38 [1837]);
assign l_37[1326]    = ( l_38 [1838]);
assign l_37[1327]    = ( l_38 [1839]);
assign l_37[1328]    = ( l_38 [1840]);
assign l_37[1329]    = ( l_38 [1841]);
assign l_37[1330]    = ( l_38 [1842]);
assign l_37[1331]    = ( l_38 [1843]);
assign l_37[1332]    = ( l_38 [1844]);
assign l_37[1333]    = ( l_38 [1845]);
assign l_37[1334]    = ( l_38 [1846]);
assign l_37[1335]    = ( l_38 [1847]);
assign l_37[1336]    = ( l_38 [1848]);
assign l_37[1337]    = ( l_38 [1849]);
assign l_37[1338]    = ( l_38 [1850]);
assign l_37[1339]    = ( l_38 [1851]);
assign l_37[1340]    = ( l_38 [1852]);
assign l_37[1341]    = ( l_38 [1853]);
assign l_37[1342]    = ( l_38 [1854]);
assign l_37[1343]    = ( l_38 [1855]);
assign l_37[1344]    = ( l_38 [1856]);
assign l_37[1345]    = ( l_38 [1857]);
assign l_37[1346]    = ( l_38 [1858]);
assign l_37[1347]    = ( l_38 [1859]);
assign l_37[1348]    = ( l_38 [1860]);
assign l_37[1349]    = ( l_38 [1861]);
assign l_37[1350]    = ( l_38 [1862]);
assign l_37[1351]    = ( l_38 [1863]);
assign l_37[1352]    = ( l_38 [1864]);
assign l_37[1353]    = ( l_38 [1865]);
assign l_37[1354]    = ( l_38 [1866]);
assign l_37[1355]    = ( l_38 [1867]);
assign l_37[1356]    = ( l_38 [1868]);
assign l_37[1357]    = ( l_38 [1869]);
assign l_37[1358]    = ( l_38 [1870]);
assign l_37[1359]    = ( l_38 [1871]);
assign l_37[1360]    = ( l_38 [1872]);
assign l_37[1361]    = ( l_38 [1873]);
assign l_37[1362]    = ( l_38 [1874]);
assign l_37[1363]    = ( l_38 [1875]);
assign l_37[1364]    = ( l_38 [1876]);
assign l_37[1365]    = ( l_38 [1877]);
assign l_37[1366]    = ( l_38 [1878]);
assign l_37[1367]    = ( l_38 [1879]);
assign l_37[1368]    = ( l_38 [1880]);
assign l_37[1369]    = ( l_38 [1881]);
assign l_37[1370]    = ( l_38 [1882]);
assign l_37[1371]    = ( l_38 [1883]);
assign l_37[1372]    = ( l_38 [1884]);
assign l_37[1373]    = ( l_38 [1885]);
assign l_37[1374]    = ( l_38 [1886]);
assign l_37[1375]    = ( l_38 [1887]);
assign l_37[1376]    = ( l_38 [1888]);
assign l_37[1377]    = ( l_38 [1889]);
assign l_37[1378]    = ( l_38 [1890]);
assign l_37[1379]    = ( l_38 [1891]);
assign l_37[1380]    = ( l_38 [1892]);
assign l_37[1381]    = ( l_38 [1893]);
assign l_37[1382]    = ( l_38 [1894]);
assign l_37[1383]    = ( l_38 [1895]);
assign l_37[1384]    = ( l_38 [1896]);
assign l_37[1385]    = ( l_38 [1897]);
assign l_37[1386]    = ( l_38 [1898]);
assign l_37[1387]    = ( l_38 [1899]);
assign l_37[1388]    = ( l_38 [1900]);
assign l_37[1389]    = ( l_38 [1901]);
assign l_37[1390]    = ( l_38 [1902]);
assign l_37[1391]    = ( l_38 [1903]);
assign l_37[1392]    = ( l_38 [1904]);
assign l_37[1393]    = ( l_38 [1905]);
assign l_37[1394]    = ( l_38 [1906]);
assign l_37[1395]    = ( l_38 [1907]);
assign l_37[1396]    = ( l_38 [1908]);
assign l_37[1397]    = ( l_38 [1909]);
assign l_37[1398]    = ( l_38 [1910]);
assign l_37[1399]    = ( l_38 [1911]);
assign l_37[1400]    = ( l_38 [1912]);
assign l_37[1401]    = ( l_38 [1913]);
assign l_37[1402]    = ( l_38 [1914]);
assign l_37[1403]    = ( l_38 [1915]);
assign l_37[1404]    = ( l_38 [1916]);
assign l_37[1405]    = ( l_38 [1917]);
assign l_37[1406]    = ( l_38 [1918]);
assign l_37[1407]    = ( l_38 [1919]);
assign l_37[1408]    = ( l_38 [1920]);
assign l_37[1409]    = ( l_38 [1921]);
assign l_37[1410]    = ( l_38 [1922]);
assign l_37[1411]    = ( l_38 [1923]);
assign l_37[1412]    = ( l_38 [1924]);
assign l_37[1413]    = ( l_38 [1925]);
assign l_37[1414]    = ( l_38 [1926]);
assign l_37[1415]    = ( l_38 [1927]);
assign l_37[1416]    = ( l_38 [1928]);
assign l_37[1417]    = ( l_38 [1929]);
assign l_37[1418]    = ( l_38 [1930]);
assign l_37[1419]    = ( l_38 [1931]);
assign l_37[1420]    = ( l_38 [1932]);
assign l_37[1421]    = ( l_38 [1933]);
assign l_37[1422]    = ( l_38 [1934]);
assign l_37[1423]    = ( l_38 [1935]);
assign l_37[1424]    = ( l_38 [1936]);
assign l_37[1425]    = ( l_38 [1937]);
assign l_37[1426]    = ( l_38 [1938]);
assign l_37[1427]    = ( l_38 [1939]);
assign l_37[1428]    = ( l_38 [1940]);
assign l_37[1429]    = ( l_38 [1941]);
assign l_37[1430]    = ( l_38 [1942]);
assign l_37[1431]    = ( l_38 [1943]);
assign l_37[1432]    = ( l_38 [1944]);
assign l_37[1433]    = ( l_38 [1945]);
assign l_37[1434]    = ( l_38 [1946]);
assign l_37[1435]    = ( l_38 [1947]);
assign l_37[1436]    = ( l_38 [1948]);
assign l_37[1437]    = ( l_38 [1949]);
assign l_37[1438]    = ( l_38 [1950]);
assign l_37[1439]    = ( l_38 [1951]);
assign l_37[1440]    = ( l_38 [1952]);
assign l_37[1441]    = ( l_38 [1953]);
assign l_37[1442]    = ( l_38 [1954]);
assign l_37[1443]    = ( l_38 [1955]);
assign l_37[1444]    = ( l_38 [1956]);
assign l_37[1445]    = ( l_38 [1957]);
assign l_37[1446]    = ( l_38 [1958]);
assign l_37[1447]    = ( l_38 [1959]);
assign l_37[1448]    = ( l_38 [1960]);
assign l_37[1449]    = ( l_38 [1961]);
assign l_37[1450]    = ( l_38 [1962]);
assign l_37[1451]    = ( l_38 [1963]);
assign l_37[1452]    = ( l_38 [1964]);
assign l_37[1453]    = ( l_38 [1965]);
assign l_37[1454]    = ( l_38 [1966]);
assign l_37[1455]    = ( l_38 [1967]);
assign l_37[1456]    = ( l_38 [1968]);
assign l_37[1457]    = ( l_38 [1969]);
assign l_37[1458]    = ( l_38 [1970]);
assign l_37[1459]    = ( l_38 [1971]);
assign l_37[1460]    = ( l_38 [1972]);
assign l_37[1461]    = ( l_38 [1973]);
assign l_37[1462]    = ( l_38 [1974]);
assign l_37[1463]    = ( l_38 [1975]);
assign l_37[1464]    = ( l_38 [1976]);
assign l_37[1465]    = ( l_38 [1977]);
assign l_37[1466]    = ( l_38 [1978]);
assign l_37[1467]    = ( l_38 [1979]);
assign l_37[1468]    = ( l_38 [1980]);
assign l_37[1469]    = ( l_38 [1981]);
assign l_37[1470]    = ( l_38 [1982]);
assign l_37[1471]    = ( l_38 [1983]);
assign l_37[1472]    = ( l_38 [1984]);
assign l_37[1473]    = ( l_38 [1985]);
assign l_37[1474]    = ( l_38 [1986]);
assign l_37[1475]    = ( l_38 [1987]);
assign l_37[1476]    = ( l_38 [1988]);
assign l_37[1477]    = ( l_38 [1989]);
assign l_37[1478]    = ( l_38 [1990]);
assign l_37[1479]    = ( l_38 [1991]);
assign l_37[1480]    = ( l_38 [1992]);
assign l_37[1481]    = ( l_38 [1993]);
assign l_37[1482]    = ( l_38 [1994]);
assign l_37[1483]    = ( l_38 [1995]);
assign l_37[1484]    = ( l_38 [1996]);
assign l_37[1485]    = ( l_38 [1997]);
assign l_37[1486]    = ( l_38 [1998]);
assign l_37[1487]    = ( l_38 [1999]);
assign l_37[1488]    = ( l_38 [2000]);
assign l_37[1489]    = ( l_38 [2001]);
assign l_37[1490]    = ( l_38 [2002]);
assign l_37[1491]    = ( l_38 [2003]);
assign l_37[1492]    = ( l_38 [2004]);
assign l_37[1493]    = ( l_38 [2005]);
assign l_37[1494]    = ( l_38 [2006]);
assign l_37[1495]    = ( l_38 [2007]);
assign l_37[1496]    = ( l_38 [2008]);
assign l_37[1497]    = ( l_38 [2009]);
assign l_37[1498]    = ( l_38 [2010]);
assign l_37[1499]    = ( l_38 [2011]);
assign l_37[1500]    = ( l_38 [2012]);
assign l_37[1501]    = ( l_38 [2013]);
assign l_37[1502]    = ( l_38 [2014]);
assign l_37[1503]    = ( l_38 [2015]);
assign l_37[1504]    = ( l_38 [2016]);
assign l_37[1505]    = ( l_38 [2017]);
assign l_37[1506]    = ( l_38 [2018]);
assign l_37[1507]    = ( l_38 [2019]);
assign l_37[1508]    = ( l_38 [2020]);
assign l_37[1509]    = ( l_38 [2021]);
assign l_37[1510]    = ( l_38 [2022]);
assign l_37[1511]    = ( l_38 [2023]);
assign l_37[1512]    = ( l_38 [2024]);
assign l_37[1513]    = ( l_38 [2025]);
assign l_37[1514]    = ( l_38 [2026]);
assign l_37[1515]    = ( l_38 [2027]);
assign l_37[1516]    = ( l_38 [2028]);
assign l_37[1517]    = ( l_38 [2029]);
assign l_37[1518]    = ( l_38 [2030]);
assign l_37[1519]    = ( l_38 [2031]);
assign l_37[1520]    = ( l_38 [2032]);
assign l_37[1521]    = ( l_38 [2033]);
assign l_37[1522]    = ( l_38 [2034]);
assign l_37[1523]    = ( l_38 [2035]);
assign l_37[1524]    = ( l_38 [2036]);
assign l_37[1525]    = ( l_38 [2037]);
assign l_37[1526]    = ( l_38 [2038]);
assign l_37[1527]    = ( l_38 [2039]);
assign l_37[1528]    = ( l_38 [2040]);
assign l_37[1529]    = ( l_38 [2041]);
assign l_37[1530]    = ( l_38 [2042]);
assign l_37[1531]    = ( l_38 [2043]);
assign l_37[1532]    = ( l_38 [2044]);
assign l_37[1533]    = ( l_38 [2045]);
assign l_37[1534]    = ( l_38 [2046]);
assign l_37[1535]    = ( l_38 [2047]);
assign l_37[1536]    = ( l_38 [2048]);
assign l_37[1537]    = ( l_38 [2049]);
assign l_37[1538]    = ( l_38 [2050]);
assign l_37[1539]    = ( l_38 [2051]);
assign l_37[1540]    = ( l_38 [2052]);
assign l_37[1541]    = ( l_38 [2053]);
assign l_37[1542]    = ( l_38 [2054]);
assign l_37[1543]    = ( l_38 [2055]);
assign l_37[1544]    = ( l_38 [2056]);
assign l_37[1545]    = ( l_38 [2057]);
assign l_37[1546]    = ( l_38 [2058]);
assign l_37[1547]    = ( l_38 [2059]);
assign l_37[1548]    = ( l_38 [2060]);
assign l_37[1549]    = ( l_38 [2061]);
assign l_37[1550]    = ( l_38 [2062]);
assign l_37[1551]    = ( l_38 [2063]);
assign l_37[1552]    = ( l_38 [2064]);
assign l_37[1553]    = ( l_38 [2065]);
assign l_38[0]    = ( l_39 [0]);
assign l_38[1]    = ( l_39 [1] & !i[1814]);
assign l_38[2]    = ( l_39 [2] & !i[1814]);
assign l_38[3]    = (!i[1814]) | ( l_39 [3] &  i[1814]);
assign l_38[4]    = (!i[1814]) | ( l_39 [4] &  i[1814]);
assign l_38[5]    = ( l_39 [5] & !i[1814]);
assign l_38[6]    = ( l_39 [6] & !i[1814]);
assign l_38[7]    = (!i[1814]) | ( l_39 [7] &  i[1814]);
assign l_38[8]    = (!i[1814]) | ( l_39 [8] &  i[1814]);
assign l_38[9]    = ( l_39 [9] & !i[1814]) | ( l_39 [10] &  i[1814]);
assign l_38[10]    = ( l_39 [10]);
assign l_38[11]    = ( l_39 [11] & !i[1814]) | ( l_39 [10] &  i[1814]);
assign l_38[12]    = ( l_39 [10] & !i[1814]) | ( l_39 [12] &  i[1814]);
assign l_38[13]    = ( l_39 [10] & !i[1814]) | ( l_39 [13] &  i[1814]);
assign l_38[14]    = ( l_39 [14] & !i[1814]) | ( l_39 [10] &  i[1814]);
assign l_38[15]    = ( l_39 [15] & !i[1814]) | ( l_39 [10] &  i[1814]);
assign l_38[16]    = ( l_39 [10] & !i[1814]) | ( l_39 [16] &  i[1814]);
assign l_38[17]    = ( l_39 [10] & !i[1814]) | ( l_39 [17] &  i[1814]);
assign l_38[18]    = ( l_39 [18]);
assign l_38[19]    = ( l_39 [19]);
assign l_38[20]    = ( l_39 [20]);
assign l_38[21]    = ( l_39 [21]);
assign l_38[22]    = ( l_39 [22]);
assign l_38[23]    = ( l_39 [23]);
assign l_38[24]    = ( l_39 [24]);
assign l_38[25]    = ( l_39 [25]);
assign l_38[26]    = ( l_39 [26]);
assign l_38[27]    = ( l_39 [27]);
assign l_38[28]    = ( l_39 [28]);
assign l_38[29]    = ( l_39 [29]);
assign l_38[30]    = ( l_39 [30]);
assign l_38[31]    = ( l_39 [31]);
assign l_38[32]    = ( l_39 [32]);
assign l_38[33]    = ( l_39 [33]);
assign l_38[34]    = ( l_39 [34]);
assign l_38[35]    = ( l_39 [35]);
assign l_38[36]    = ( l_39 [36]);
assign l_38[37]    = ( l_39 [37]);
assign l_38[38]    = ( l_39 [38]);
assign l_38[39]    = ( l_39 [39]);
assign l_38[40]    = ( l_39 [40]);
assign l_38[41]    = ( l_39 [41]);
assign l_38[42]    = ( l_39 [42]);
assign l_38[43]    = ( l_39 [43]);
assign l_38[44]    = ( l_39 [44]);
assign l_38[45]    = ( l_39 [45]);
assign l_38[46]    = ( l_39 [46]);
assign l_38[47]    = ( l_39 [47]);
assign l_38[48]    = ( l_39 [48]);
assign l_38[49]    = ( l_39 [49]);
assign l_38[50]    = ( l_39 [50]);
assign l_38[51]    = ( l_39 [51]);
assign l_38[52]    = ( l_39 [52]);
assign l_38[53]    = ( l_39 [53]);
assign l_38[54]    = ( l_39 [54]);
assign l_38[55]    = ( l_39 [55]);
assign l_38[56]    = ( l_39 [56]);
assign l_38[57]    = ( l_39 [57]);
assign l_38[58]    = ( l_39 [58]);
assign l_38[59]    = ( l_39 [59]);
assign l_38[60]    = ( l_39 [60]);
assign l_38[61]    = ( l_39 [61]);
assign l_38[62]    = ( l_39 [62]);
assign l_38[63]    = ( l_39 [63]);
assign l_38[64]    = ( l_39 [64]);
assign l_38[65]    = ( l_39 [65]);
assign l_38[66]    = ( l_39 [66]);
assign l_38[67]    = ( l_39 [67]);
assign l_38[68]    = ( l_39 [68]);
assign l_38[69]    = ( l_39 [69]);
assign l_38[70]    = ( l_39 [70]);
assign l_38[71]    = ( l_39 [71]);
assign l_38[72]    = ( l_39 [72]);
assign l_38[73]    = ( l_39 [73]);
assign l_38[74]    = ( l_39 [74]);
assign l_38[75]    = ( l_39 [75]);
assign l_38[76]    = ( l_39 [76]);
assign l_38[77]    = ( l_39 [77]);
assign l_38[78]    = ( l_39 [78]);
assign l_38[79]    = ( l_39 [79]);
assign l_38[80]    = ( l_39 [80]);
assign l_38[81]    = ( l_39 [81]);
assign l_38[82]    = ( l_39 [82]);
assign l_38[83]    = ( l_39 [83]);
assign l_38[84]    = ( l_39 [84]);
assign l_38[85]    = ( l_39 [85]);
assign l_38[86]    = ( l_39 [86]);
assign l_38[87]    = ( l_39 [87]);
assign l_38[88]    = ( l_39 [88]);
assign l_38[89]    = ( l_39 [89]);
assign l_38[90]    = ( l_39 [90]);
assign l_38[91]    = ( l_39 [91]);
assign l_38[92]    = ( l_39 [92]);
assign l_38[93]    = ( l_39 [93]);
assign l_38[94]    = ( l_39 [94]);
assign l_38[95]    = ( l_39 [95]);
assign l_38[96]    = ( l_39 [96]);
assign l_38[97]    = ( l_39 [97]);
assign l_38[98]    = ( l_39 [98]);
assign l_38[99]    = ( l_39 [99]);
assign l_38[100]    = ( l_39 [100]);
assign l_38[101]    = ( l_39 [101]);
assign l_38[102]    = ( l_39 [102]);
assign l_38[103]    = ( l_39 [103]);
assign l_38[104]    = ( l_39 [104]);
assign l_38[105]    = ( l_39 [105]);
assign l_38[106]    = ( l_39 [106]);
assign l_38[107]    = ( l_39 [107]);
assign l_38[108]    = ( l_39 [108]);
assign l_38[109]    = ( l_39 [109]);
assign l_38[110]    = ( l_39 [110]);
assign l_38[111]    = ( l_39 [111]);
assign l_38[112]    = ( l_39 [112]);
assign l_38[113]    = ( l_39 [113]);
assign l_38[114]    = ( l_39 [114]);
assign l_38[115]    = ( l_39 [115]);
assign l_38[116]    = ( l_39 [116]);
assign l_38[117]    = ( l_39 [117]);
assign l_38[118]    = ( l_39 [118]);
assign l_38[119]    = ( l_39 [119]);
assign l_38[120]    = ( l_39 [120]);
assign l_38[121]    = ( l_39 [121]);
assign l_38[122]    = ( l_39 [122]);
assign l_38[123]    = ( l_39 [123]);
assign l_38[124]    = ( l_39 [124]);
assign l_38[125]    = ( l_39 [125]);
assign l_38[126]    = ( l_39 [126]);
assign l_38[127]    = ( l_39 [127]);
assign l_38[128]    = ( l_39 [128]);
assign l_38[129]    = ( l_39 [129]);
assign l_38[130]    = ( l_39 [130]);
assign l_38[131]    = ( l_39 [131]);
assign l_38[132]    = ( l_39 [132]);
assign l_38[133]    = ( l_39 [133]);
assign l_38[134]    = ( l_39 [134]);
assign l_38[135]    = ( l_39 [135]);
assign l_38[136]    = ( l_39 [136]);
assign l_38[137]    = ( l_39 [137]);
assign l_38[138]    = ( l_39 [138]);
assign l_38[139]    = ( l_39 [139]);
assign l_38[140]    = ( l_39 [140]);
assign l_38[141]    = ( l_39 [141]);
assign l_38[142]    = ( l_39 [142]);
assign l_38[143]    = ( l_39 [143]);
assign l_38[144]    = ( l_39 [144]);
assign l_38[145]    = ( l_39 [145]);
assign l_38[146]    = ( l_39 [146]);
assign l_38[147]    = ( l_39 [147]);
assign l_38[148]    = ( l_39 [148]);
assign l_38[149]    = ( l_39 [149]);
assign l_38[150]    = ( l_39 [150]);
assign l_38[151]    = ( l_39 [151]);
assign l_38[152]    = ( l_39 [152]);
assign l_38[153]    = ( l_39 [153]);
assign l_38[154]    = ( l_39 [154]);
assign l_38[155]    = ( l_39 [155]);
assign l_38[156]    = ( l_39 [156]);
assign l_38[157]    = ( l_39 [157]);
assign l_38[158]    = ( l_39 [158]);
assign l_38[159]    = ( l_39 [159]);
assign l_38[160]    = ( l_39 [160]);
assign l_38[161]    = ( l_39 [161]);
assign l_38[162]    = ( l_39 [162]);
assign l_38[163]    = ( l_39 [163]);
assign l_38[164]    = ( l_39 [164]);
assign l_38[165]    = ( l_39 [165]);
assign l_38[166]    = ( l_39 [166]);
assign l_38[167]    = ( l_39 [167]);
assign l_38[168]    = ( l_39 [168]);
assign l_38[169]    = ( l_39 [169]);
assign l_38[170]    = ( l_39 [170]);
assign l_38[171]    = ( l_39 [171]);
assign l_38[172]    = ( l_39 [172]);
assign l_38[173]    = ( l_39 [173]);
assign l_38[174]    = ( l_39 [174]);
assign l_38[175]    = ( l_39 [175]);
assign l_38[176]    = ( l_39 [176]);
assign l_38[177]    = ( l_39 [177]);
assign l_38[178]    = ( l_39 [178]);
assign l_38[179]    = ( l_39 [179]);
assign l_38[180]    = ( l_39 [180]);
assign l_38[181]    = ( l_39 [181]);
assign l_38[182]    = ( l_39 [182]);
assign l_38[183]    = ( l_39 [183]);
assign l_38[184]    = ( l_39 [184]);
assign l_38[185]    = ( l_39 [185]);
assign l_38[186]    = ( l_39 [186]);
assign l_38[187]    = ( l_39 [187]);
assign l_38[188]    = ( l_39 [188]);
assign l_38[189]    = ( l_39 [189]);
assign l_38[190]    = ( l_39 [190]);
assign l_38[191]    = ( l_39 [191]);
assign l_38[192]    = ( l_39 [192]);
assign l_38[193]    = ( l_39 [193]);
assign l_38[194]    = ( l_39 [194]);
assign l_38[195]    = ( l_39 [195]);
assign l_38[196]    = ( l_39 [196]);
assign l_38[197]    = ( l_39 [197]);
assign l_38[198]    = ( l_39 [198]);
assign l_38[199]    = ( l_39 [199]);
assign l_38[200]    = ( l_39 [200]);
assign l_38[201]    = ( l_39 [201]);
assign l_38[202]    = ( l_39 [202]);
assign l_38[203]    = ( l_39 [203]);
assign l_38[204]    = ( l_39 [204]);
assign l_38[205]    = ( l_39 [205]);
assign l_38[206]    = ( l_39 [206]);
assign l_38[207]    = ( l_39 [207]);
assign l_38[208]    = ( l_39 [208]);
assign l_38[209]    = ( l_39 [209]);
assign l_38[210]    = ( l_39 [210]);
assign l_38[211]    = ( l_39 [211]);
assign l_38[212]    = ( l_39 [212]);
assign l_38[213]    = ( l_39 [213]);
assign l_38[214]    = ( l_39 [214]);
assign l_38[215]    = ( l_39 [215]);
assign l_38[216]    = ( l_39 [216]);
assign l_38[217]    = ( l_39 [217]);
assign l_38[218]    = ( l_39 [218]);
assign l_38[219]    = ( l_39 [219]);
assign l_38[220]    = ( l_39 [220]);
assign l_38[221]    = ( l_39 [221]);
assign l_38[222]    = ( l_39 [222]);
assign l_38[223]    = ( l_39 [223]);
assign l_38[224]    = ( l_39 [224]);
assign l_38[225]    = ( l_39 [225]);
assign l_38[226]    = ( l_39 [226]);
assign l_38[227]    = ( l_39 [227]);
assign l_38[228]    = ( l_39 [228]);
assign l_38[229]    = ( l_39 [229]);
assign l_38[230]    = ( l_39 [230]);
assign l_38[231]    = ( l_39 [231]);
assign l_38[232]    = ( l_39 [232]);
assign l_38[233]    = ( l_39 [233]);
assign l_38[234]    = ( l_39 [234]);
assign l_38[235]    = ( l_39 [235]);
assign l_38[236]    = ( l_39 [236]);
assign l_38[237]    = ( l_39 [237]);
assign l_38[238]    = ( l_39 [238]);
assign l_38[239]    = ( l_39 [239]);
assign l_38[240]    = ( l_39 [240]);
assign l_38[241]    = ( l_39 [241]);
assign l_38[242]    = ( l_39 [242]);
assign l_38[243]    = ( l_39 [243]);
assign l_38[244]    = ( l_39 [244]);
assign l_38[245]    = ( l_39 [245]);
assign l_38[246]    = ( l_39 [246]);
assign l_38[247]    = ( l_39 [247]);
assign l_38[248]    = ( l_39 [248]);
assign l_38[249]    = ( l_39 [249]);
assign l_38[250]    = ( l_39 [250]);
assign l_38[251]    = ( l_39 [251]);
assign l_38[252]    = ( l_39 [252]);
assign l_38[253]    = ( l_39 [253]);
assign l_38[254]    = ( l_39 [254]);
assign l_38[255]    = ( l_39 [255]);
assign l_38[256]    = ( l_39 [256]);
assign l_38[257]    = ( l_39 [257]);
assign l_38[258]    = ( l_39 [258]);
assign l_38[259]    = ( l_39 [259]);
assign l_38[260]    = ( l_39 [260]);
assign l_38[261]    = ( l_39 [261]);
assign l_38[262]    = ( l_39 [262]);
assign l_38[263]    = ( l_39 [263]);
assign l_38[264]    = ( l_39 [264]);
assign l_38[265]    = ( l_39 [265]);
assign l_38[266]    = ( l_39 [266]);
assign l_38[267]    = ( l_39 [267]);
assign l_38[268]    = ( l_39 [268]);
assign l_38[269]    = ( l_39 [269]);
assign l_38[270]    = ( l_39 [270]);
assign l_38[271]    = ( l_39 [271]);
assign l_38[272]    = ( l_39 [272]);
assign l_38[273]    = ( l_39 [273]);
assign l_38[274]    = ( l_39 [274]);
assign l_38[275]    = ( l_39 [275]);
assign l_38[276]    = ( l_39 [276]);
assign l_38[277]    = ( l_39 [277]);
assign l_38[278]    = ( l_39 [278]);
assign l_38[279]    = ( l_39 [279]);
assign l_38[280]    = ( l_39 [280]);
assign l_38[281]    = ( l_39 [281]);
assign l_38[282]    = ( l_39 [282]);
assign l_38[283]    = ( l_39 [283]);
assign l_38[284]    = ( l_39 [284]);
assign l_38[285]    = ( l_39 [285]);
assign l_38[286]    = ( l_39 [286]);
assign l_38[287]    = ( l_39 [287]);
assign l_38[288]    = ( l_39 [288]);
assign l_38[289]    = ( l_39 [289]);
assign l_38[290]    = ( l_39 [290]);
assign l_38[291]    = ( l_39 [291]);
assign l_38[292]    = ( l_39 [292]);
assign l_38[293]    = ( l_39 [293]);
assign l_38[294]    = ( l_39 [294]);
assign l_38[295]    = ( l_39 [295]);
assign l_38[296]    = ( l_39 [296]);
assign l_38[297]    = ( l_39 [297]);
assign l_38[298]    = ( l_39 [298]);
assign l_38[299]    = ( l_39 [299]);
assign l_38[300]    = ( l_39 [300]);
assign l_38[301]    = ( l_39 [301]);
assign l_38[302]    = ( l_39 [302]);
assign l_38[303]    = ( l_39 [303]);
assign l_38[304]    = ( l_39 [304]);
assign l_38[305]    = ( l_39 [305]);
assign l_38[306]    = ( l_39 [306]);
assign l_38[307]    = ( l_39 [307]);
assign l_38[308]    = ( l_39 [308]);
assign l_38[309]    = ( l_39 [309]);
assign l_38[310]    = ( l_39 [310]);
assign l_38[311]    = ( l_39 [311]);
assign l_38[312]    = ( l_39 [312]);
assign l_38[313]    = ( l_39 [313]);
assign l_38[314]    = ( l_39 [314]);
assign l_38[315]    = ( l_39 [315]);
assign l_38[316]    = ( l_39 [316]);
assign l_38[317]    = ( l_39 [317]);
assign l_38[318]    = ( l_39 [318]);
assign l_38[319]    = ( l_39 [319]);
assign l_38[320]    = ( l_39 [320]);
assign l_38[321]    = ( l_39 [321]);
assign l_38[322]    = ( l_39 [322]);
assign l_38[323]    = ( l_39 [323]);
assign l_38[324]    = ( l_39 [324]);
assign l_38[325]    = ( l_39 [325]);
assign l_38[326]    = ( l_39 [326]);
assign l_38[327]    = ( l_39 [327]);
assign l_38[328]    = ( l_39 [328]);
assign l_38[329]    = ( l_39 [329]);
assign l_38[330]    = ( l_39 [330]);
assign l_38[331]    = ( l_39 [331]);
assign l_38[332]    = ( l_39 [332]);
assign l_38[333]    = ( l_39 [333]);
assign l_38[334]    = ( l_39 [334]);
assign l_38[335]    = ( l_39 [335]);
assign l_38[336]    = ( l_39 [336]);
assign l_38[337]    = ( l_39 [337]);
assign l_38[338]    = ( l_39 [338]);
assign l_38[339]    = ( l_39 [339]);
assign l_38[340]    = ( l_39 [340]);
assign l_38[341]    = ( l_39 [341]);
assign l_38[342]    = ( l_39 [342]);
assign l_38[343]    = ( l_39 [343]);
assign l_38[344]    = ( l_39 [344]);
assign l_38[345]    = ( l_39 [345]);
assign l_38[346]    = ( l_39 [346]);
assign l_38[347]    = ( l_39 [347]);
assign l_38[348]    = ( l_39 [348]);
assign l_38[349]    = ( l_39 [349]);
assign l_38[350]    = ( l_39 [350]);
assign l_38[351]    = ( l_39 [351]);
assign l_38[352]    = ( l_39 [352]);
assign l_38[353]    = ( l_39 [353]);
assign l_38[354]    = ( l_39 [354]);
assign l_38[355]    = ( l_39 [355]);
assign l_38[356]    = ( l_39 [356]);
assign l_38[357]    = ( l_39 [357]);
assign l_38[358]    = ( l_39 [358]);
assign l_38[359]    = ( l_39 [359]);
assign l_38[360]    = ( l_39 [360]);
assign l_38[361]    = ( l_39 [361]);
assign l_38[362]    = ( l_39 [362]);
assign l_38[363]    = ( l_39 [363]);
assign l_38[364]    = ( l_39 [364]);
assign l_38[365]    = ( l_39 [365]);
assign l_38[366]    = ( l_39 [366]);
assign l_38[367]    = ( l_39 [367]);
assign l_38[368]    = ( l_39 [368]);
assign l_38[369]    = ( l_39 [369]);
assign l_38[370]    = ( l_39 [370]);
assign l_38[371]    = ( l_39 [371]);
assign l_38[372]    = ( l_39 [372]);
assign l_38[373]    = ( l_39 [373]);
assign l_38[374]    = ( l_39 [374]);
assign l_38[375]    = ( l_39 [375]);
assign l_38[376]    = ( l_39 [376]);
assign l_38[377]    = ( l_39 [377]);
assign l_38[378]    = ( l_39 [378]);
assign l_38[379]    = ( l_39 [379]);
assign l_38[380]    = ( l_39 [380]);
assign l_38[381]    = ( l_39 [381]);
assign l_38[382]    = ( l_39 [382]);
assign l_38[383]    = ( l_39 [383]);
assign l_38[384]    = ( l_39 [384]);
assign l_38[385]    = ( l_39 [385]);
assign l_38[386]    = ( l_39 [386]);
assign l_38[387]    = ( l_39 [387]);
assign l_38[388]    = ( l_39 [388]);
assign l_38[389]    = ( l_39 [389]);
assign l_38[390]    = ( l_39 [390]);
assign l_38[391]    = ( l_39 [391]);
assign l_38[392]    = ( l_39 [392]);
assign l_38[393]    = ( l_39 [393]);
assign l_38[394]    = ( l_39 [394]);
assign l_38[395]    = ( l_39 [395]);
assign l_38[396]    = ( l_39 [396]);
assign l_38[397]    = ( l_39 [397]);
assign l_38[398]    = ( l_39 [398]);
assign l_38[399]    = ( l_39 [399]);
assign l_38[400]    = ( l_39 [400]);
assign l_38[401]    = ( l_39 [401]);
assign l_38[402]    = ( l_39 [402]);
assign l_38[403]    = ( l_39 [403]);
assign l_38[404]    = ( l_39 [404]);
assign l_38[405]    = ( l_39 [405]);
assign l_38[406]    = ( l_39 [406]);
assign l_38[407]    = ( l_39 [407]);
assign l_38[408]    = ( l_39 [408]);
assign l_38[409]    = ( l_39 [409]);
assign l_38[410]    = ( l_39 [410]);
assign l_38[411]    = ( l_39 [411]);
assign l_38[412]    = ( l_39 [412]);
assign l_38[413]    = ( l_39 [413]);
assign l_38[414]    = ( l_39 [414]);
assign l_38[415]    = ( l_39 [415]);
assign l_38[416]    = ( l_39 [416]);
assign l_38[417]    = ( l_39 [417]);
assign l_38[418]    = ( l_39 [418]);
assign l_38[419]    = ( l_39 [419]);
assign l_38[420]    = ( l_39 [420]);
assign l_38[421]    = ( l_39 [421]);
assign l_38[422]    = ( l_39 [422]);
assign l_38[423]    = ( l_39 [423]);
assign l_38[424]    = ( l_39 [424]);
assign l_38[425]    = ( l_39 [425]);
assign l_38[426]    = ( l_39 [426]);
assign l_38[427]    = ( l_39 [427]);
assign l_38[428]    = ( l_39 [428]);
assign l_38[429]    = ( l_39 [429]);
assign l_38[430]    = ( l_39 [430]);
assign l_38[431]    = ( l_39 [431]);
assign l_38[432]    = ( l_39 [432]);
assign l_38[433]    = ( l_39 [433]);
assign l_38[434]    = ( l_39 [434]);
assign l_38[435]    = ( l_39 [435]);
assign l_38[436]    = ( l_39 [436]);
assign l_38[437]    = ( l_39 [437]);
assign l_38[438]    = ( l_39 [438]);
assign l_38[439]    = ( l_39 [439]);
assign l_38[440]    = ( l_39 [440]);
assign l_38[441]    = ( l_39 [441]);
assign l_38[442]    = ( l_39 [442]);
assign l_38[443]    = ( l_39 [443]);
assign l_38[444]    = ( l_39 [444]);
assign l_38[445]    = ( l_39 [445]);
assign l_38[446]    = ( l_39 [446]);
assign l_38[447]    = ( l_39 [447]);
assign l_38[448]    = ( l_39 [448]);
assign l_38[449]    = ( l_39 [449]);
assign l_38[450]    = ( l_39 [450]);
assign l_38[451]    = ( l_39 [451]);
assign l_38[452]    = ( l_39 [452]);
assign l_38[453]    = ( l_39 [453]);
assign l_38[454]    = ( l_39 [454]);
assign l_38[455]    = ( l_39 [455]);
assign l_38[456]    = ( l_39 [456]);
assign l_38[457]    = ( l_39 [457]);
assign l_38[458]    = ( l_39 [458]);
assign l_38[459]    = ( l_39 [459]);
assign l_38[460]    = ( l_39 [460]);
assign l_38[461]    = ( l_39 [461]);
assign l_38[462]    = ( l_39 [462]);
assign l_38[463]    = ( l_39 [463]);
assign l_38[464]    = ( l_39 [464]);
assign l_38[465]    = ( l_39 [465]);
assign l_38[466]    = ( l_39 [466]);
assign l_38[467]    = ( l_39 [467]);
assign l_38[468]    = ( l_39 [468]);
assign l_38[469]    = ( l_39 [469]);
assign l_38[470]    = ( l_39 [470]);
assign l_38[471]    = ( l_39 [471]);
assign l_38[472]    = ( l_39 [472]);
assign l_38[473]    = ( l_39 [473]);
assign l_38[474]    = ( l_39 [474]);
assign l_38[475]    = ( l_39 [475]);
assign l_38[476]    = ( l_39 [476]);
assign l_38[477]    = ( l_39 [477]);
assign l_38[478]    = ( l_39 [478]);
assign l_38[479]    = ( l_39 [479]);
assign l_38[480]    = ( l_39 [480]);
assign l_38[481]    = ( l_39 [481]);
assign l_38[482]    = ( l_39 [482]);
assign l_38[483]    = ( l_39 [483]);
assign l_38[484]    = ( l_39 [484]);
assign l_38[485]    = ( l_39 [485]);
assign l_38[486]    = ( l_39 [486]);
assign l_38[487]    = ( l_39 [487]);
assign l_38[488]    = ( l_39 [488]);
assign l_38[489]    = ( l_39 [489]);
assign l_38[490]    = ( l_39 [490]);
assign l_38[491]    = ( l_39 [491]);
assign l_38[492]    = ( l_39 [492]);
assign l_38[493]    = ( l_39 [493]);
assign l_38[494]    = ( l_39 [494]);
assign l_38[495]    = ( l_39 [495]);
assign l_38[496]    = ( l_39 [496]);
assign l_38[497]    = ( l_39 [497]);
assign l_38[498]    = ( l_39 [498]);
assign l_38[499]    = ( l_39 [499]);
assign l_38[500]    = ( l_39 [500]);
assign l_38[501]    = ( l_39 [501]);
assign l_38[502]    = ( l_39 [502]);
assign l_38[503]    = ( l_39 [503]);
assign l_38[504]    = ( l_39 [504]);
assign l_38[505]    = ( l_39 [505]);
assign l_38[506]    = ( l_39 [506]);
assign l_38[507]    = ( l_39 [507]);
assign l_38[508]    = ( l_39 [508]);
assign l_38[509]    = ( l_39 [509]);
assign l_38[510]    = ( l_39 [510]);
assign l_38[511]    = ( l_39 [511]);
assign l_38[512]    = ( l_39 [512]);
assign l_38[513]    = ( l_39 [513]);
assign l_38[514]    = ( l_39 [514]);
assign l_38[515]    = ( l_39 [515]);
assign l_38[516]    = ( l_39 [516]);
assign l_38[517]    = ( l_39 [517]);
assign l_38[518]    = ( l_39 [518]);
assign l_38[519]    = ( l_39 [519]);
assign l_38[520]    = ( l_39 [520]);
assign l_38[521]    = ( l_39 [521]);
assign l_38[522]    = ( l_39 [522]);
assign l_38[523]    = ( l_39 [523]);
assign l_38[524]    = ( l_39 [524]);
assign l_38[525]    = ( l_39 [525]);
assign l_38[526]    = ( l_39 [526]);
assign l_38[527]    = ( l_39 [527]);
assign l_38[528]    = ( l_39 [528]);
assign l_38[529]    = ( l_39 [529]);
assign l_38[530]    = ( l_39 [530]);
assign l_38[531]    = ( l_39 [531]);
assign l_38[532]    = ( l_39 [532]);
assign l_38[533]    = ( l_39 [533]);
assign l_38[534]    = ( l_39 [534]);
assign l_38[535]    = ( l_39 [535]);
assign l_38[536]    = ( l_39 [536]);
assign l_38[537]    = ( l_39 [537]);
assign l_38[538]    = ( l_39 [538]);
assign l_38[539]    = ( l_39 [539]);
assign l_38[540]    = ( l_39 [540]);
assign l_38[541]    = ( l_39 [541]);
assign l_38[542]    = ( l_39 [542]);
assign l_38[543]    = ( l_39 [543]);
assign l_38[544]    = ( l_39 [544]);
assign l_38[545]    = ( l_39 [545]);
assign l_38[546]    = ( l_39 [546]);
assign l_38[547]    = ( l_39 [547]);
assign l_38[548]    = ( l_39 [548]);
assign l_38[549]    = ( l_39 [549]);
assign l_38[550]    = ( l_39 [550]);
assign l_38[551]    = ( l_39 [551]);
assign l_38[552]    = ( l_39 [552]);
assign l_38[553]    = ( l_39 [553]);
assign l_38[554]    = ( l_39 [554]);
assign l_38[555]    = ( l_39 [555]);
assign l_38[556]    = ( l_39 [556]);
assign l_38[557]    = ( l_39 [557]);
assign l_38[558]    = ( l_39 [558]);
assign l_38[559]    = ( l_39 [559]);
assign l_38[560]    = ( l_39 [560]);
assign l_38[561]    = ( l_39 [561]);
assign l_38[562]    = ( l_39 [562]);
assign l_38[563]    = ( l_39 [563]);
assign l_38[564]    = ( l_39 [564]);
assign l_38[565]    = ( l_39 [565]);
assign l_38[566]    = ( l_39 [566]);
assign l_38[567]    = ( l_39 [567]);
assign l_38[568]    = ( l_39 [568]);
assign l_38[569]    = ( l_39 [569]);
assign l_38[570]    = ( l_39 [570]);
assign l_38[571]    = ( l_39 [571]);
assign l_38[572]    = ( l_39 [572]);
assign l_38[573]    = ( l_39 [573]);
assign l_38[574]    = ( l_39 [574]);
assign l_38[575]    = ( l_39 [575]);
assign l_38[576]    = ( l_39 [576]);
assign l_38[577]    = ( l_39 [577]);
assign l_38[578]    = ( l_39 [578]);
assign l_38[579]    = ( l_39 [579]);
assign l_38[580]    = ( l_39 [580]);
assign l_38[581]    = ( l_39 [581]);
assign l_38[582]    = ( l_39 [582]);
assign l_38[583]    = ( l_39 [583]);
assign l_38[584]    = ( l_39 [584]);
assign l_38[585]    = ( l_39 [585]);
assign l_38[586]    = ( l_39 [586]);
assign l_38[587]    = ( l_39 [587]);
assign l_38[588]    = ( l_39 [588]);
assign l_38[589]    = ( l_39 [589]);
assign l_38[590]    = ( l_39 [590]);
assign l_38[591]    = ( l_39 [591]);
assign l_38[592]    = ( l_39 [592]);
assign l_38[593]    = ( l_39 [593]);
assign l_38[594]    = ( l_39 [594]);
assign l_38[595]    = ( l_39 [595]);
assign l_38[596]    = ( l_39 [596]);
assign l_38[597]    = ( l_39 [597]);
assign l_38[598]    = ( l_39 [598]);
assign l_38[599]    = ( l_39 [599]);
assign l_38[600]    = ( l_39 [600]);
assign l_38[601]    = ( l_39 [601]);
assign l_38[602]    = ( l_39 [602]);
assign l_38[603]    = ( l_39 [603]);
assign l_38[604]    = ( l_39 [604]);
assign l_38[605]    = ( l_39 [605]);
assign l_38[606]    = ( l_39 [606]);
assign l_38[607]    = ( l_39 [607]);
assign l_38[608]    = ( l_39 [608]);
assign l_38[609]    = ( l_39 [609]);
assign l_38[610]    = ( l_39 [610]);
assign l_38[611]    = ( l_39 [611]);
assign l_38[612]    = ( l_39 [612]);
assign l_38[613]    = ( l_39 [613]);
assign l_38[614]    = ( l_39 [614]);
assign l_38[615]    = ( l_39 [615]);
assign l_38[616]    = ( l_39 [616]);
assign l_38[617]    = ( l_39 [617]);
assign l_38[618]    = ( l_39 [618]);
assign l_38[619]    = ( l_39 [619]);
assign l_38[620]    = ( l_39 [620]);
assign l_38[621]    = ( l_39 [621]);
assign l_38[622]    = ( l_39 [622]);
assign l_38[623]    = ( l_39 [623]);
assign l_38[624]    = ( l_39 [624]);
assign l_38[625]    = ( l_39 [625]);
assign l_38[626]    = ( l_39 [626]);
assign l_38[627]    = ( l_39 [627]);
assign l_38[628]    = ( l_39 [628]);
assign l_38[629]    = ( l_39 [629]);
assign l_38[630]    = ( l_39 [630]);
assign l_38[631]    = ( l_39 [631]);
assign l_38[632]    = ( l_39 [632]);
assign l_38[633]    = ( l_39 [633]);
assign l_38[634]    = ( l_39 [634]);
assign l_38[635]    = ( l_39 [635]);
assign l_38[636]    = ( l_39 [636]);
assign l_38[637]    = ( l_39 [637]);
assign l_38[638]    = ( l_39 [638]);
assign l_38[639]    = ( l_39 [639]);
assign l_38[640]    = ( l_39 [640]);
assign l_38[641]    = ( l_39 [641]);
assign l_38[642]    = ( l_39 [642]);
assign l_38[643]    = ( l_39 [643]);
assign l_38[644]    = ( l_39 [644]);
assign l_38[645]    = ( l_39 [645]);
assign l_38[646]    = ( l_39 [646]);
assign l_38[647]    = ( l_39 [647]);
assign l_38[648]    = ( l_39 [648]);
assign l_38[649]    = ( l_39 [649]);
assign l_38[650]    = ( l_39 [650]);
assign l_38[651]    = ( l_39 [651]);
assign l_38[652]    = ( l_39 [652]);
assign l_38[653]    = ( l_39 [653]);
assign l_38[654]    = ( l_39 [654]);
assign l_38[655]    = ( l_39 [655]);
assign l_38[656]    = ( l_39 [656]);
assign l_38[657]    = ( l_39 [657]);
assign l_38[658]    = ( l_39 [658]);
assign l_38[659]    = ( l_39 [659]);
assign l_38[660]    = ( l_39 [660]);
assign l_38[661]    = ( l_39 [661]);
assign l_38[662]    = ( l_39 [662]);
assign l_38[663]    = ( l_39 [663]);
assign l_38[664]    = ( l_39 [664]);
assign l_38[665]    = ( l_39 [665]);
assign l_38[666]    = ( l_39 [666]);
assign l_38[667]    = ( l_39 [667]);
assign l_38[668]    = ( l_39 [668]);
assign l_38[669]    = ( l_39 [669]);
assign l_38[670]    = ( l_39 [670]);
assign l_38[671]    = ( l_39 [671]);
assign l_38[672]    = ( l_39 [672]);
assign l_38[673]    = ( l_39 [673]);
assign l_38[674]    = ( l_39 [674]);
assign l_38[675]    = ( l_39 [675]);
assign l_38[676]    = ( l_39 [676]);
assign l_38[677]    = ( l_39 [677]);
assign l_38[678]    = ( l_39 [678]);
assign l_38[679]    = ( l_39 [679]);
assign l_38[680]    = ( l_39 [680]);
assign l_38[681]    = ( l_39 [681]);
assign l_38[682]    = ( l_39 [682]);
assign l_38[683]    = ( l_39 [683]);
assign l_38[684]    = ( l_39 [684]);
assign l_38[685]    = ( l_39 [685]);
assign l_38[686]    = ( l_39 [686]);
assign l_38[687]    = ( l_39 [687]);
assign l_38[688]    = ( l_39 [688]);
assign l_38[689]    = ( l_39 [689]);
assign l_38[690]    = ( l_39 [690]);
assign l_38[691]    = ( l_39 [691]);
assign l_38[692]    = ( l_39 [692]);
assign l_38[693]    = ( l_39 [693]);
assign l_38[694]    = ( l_39 [694]);
assign l_38[695]    = ( l_39 [695]);
assign l_38[696]    = ( l_39 [696]);
assign l_38[697]    = ( l_39 [697]);
assign l_38[698]    = ( l_39 [698]);
assign l_38[699]    = ( l_39 [699]);
assign l_38[700]    = ( l_39 [700]);
assign l_38[701]    = ( l_39 [701]);
assign l_38[702]    = ( l_39 [702]);
assign l_38[703]    = ( l_39 [703]);
assign l_38[704]    = ( l_39 [704]);
assign l_38[705]    = ( l_39 [705]);
assign l_38[706]    = ( l_39 [706]);
assign l_38[707]    = ( l_39 [707]);
assign l_38[708]    = ( l_39 [708]);
assign l_38[709]    = ( l_39 [709]);
assign l_38[710]    = ( l_39 [710]);
assign l_38[711]    = ( l_39 [711]);
assign l_38[712]    = ( l_39 [712]);
assign l_38[713]    = ( l_39 [713]);
assign l_38[714]    = ( l_39 [714]);
assign l_38[715]    = ( l_39 [715]);
assign l_38[716]    = ( l_39 [716]);
assign l_38[717]    = ( l_39 [717]);
assign l_38[718]    = ( l_39 [718]);
assign l_38[719]    = ( l_39 [719]);
assign l_38[720]    = ( l_39 [720]);
assign l_38[721]    = ( l_39 [721]);
assign l_38[722]    = ( l_39 [722]);
assign l_38[723]    = ( l_39 [723]);
assign l_38[724]    = ( l_39 [724]);
assign l_38[725]    = ( l_39 [725]);
assign l_38[726]    = ( l_39 [726]);
assign l_38[727]    = ( l_39 [727]);
assign l_38[728]    = ( l_39 [728]);
assign l_38[729]    = ( l_39 [729]);
assign l_38[730]    = ( l_39 [730]);
assign l_38[731]    = ( l_39 [731]);
assign l_38[732]    = ( l_39 [732]);
assign l_38[733]    = ( l_39 [733]);
assign l_38[734]    = ( l_39 [734]);
assign l_38[735]    = ( l_39 [735]);
assign l_38[736]    = ( l_39 [736]);
assign l_38[737]    = ( l_39 [737]);
assign l_38[738]    = ( l_39 [738]);
assign l_38[739]    = ( l_39 [739]);
assign l_38[740]    = ( l_39 [740]);
assign l_38[741]    = ( l_39 [741]);
assign l_38[742]    = ( l_39 [742]);
assign l_38[743]    = ( l_39 [743]);
assign l_38[744]    = ( l_39 [744]);
assign l_38[745]    = ( l_39 [745]);
assign l_38[746]    = ( l_39 [746]);
assign l_38[747]    = ( l_39 [747]);
assign l_38[748]    = ( l_39 [748]);
assign l_38[749]    = ( l_39 [749]);
assign l_38[750]    = ( l_39 [750]);
assign l_38[751]    = ( l_39 [751]);
assign l_38[752]    = ( l_39 [752]);
assign l_38[753]    = ( l_39 [753]);
assign l_38[754]    = ( l_39 [754]);
assign l_38[755]    = ( l_39 [755]);
assign l_38[756]    = ( l_39 [756]);
assign l_38[757]    = ( l_39 [757]);
assign l_38[758]    = ( l_39 [758]);
assign l_38[759]    = ( l_39 [759]);
assign l_38[760]    = ( l_39 [760]);
assign l_38[761]    = ( l_39 [761]);
assign l_38[762]    = ( l_39 [762]);
assign l_38[763]    = ( l_39 [763]);
assign l_38[764]    = ( l_39 [764]);
assign l_38[765]    = ( l_39 [765]);
assign l_38[766]    = ( l_39 [766]);
assign l_38[767]    = ( l_39 [767]);
assign l_38[768]    = ( l_39 [768]);
assign l_38[769]    = ( l_39 [769]);
assign l_38[770]    = ( l_39 [770]);
assign l_38[771]    = ( l_39 [771]);
assign l_38[772]    = ( l_39 [772]);
assign l_38[773]    = ( l_39 [773]);
assign l_38[774]    = ( l_39 [774]);
assign l_38[775]    = ( l_39 [775]);
assign l_38[776]    = ( l_39 [776]);
assign l_38[777]    = ( l_39 [777]);
assign l_38[778]    = ( l_39 [778]);
assign l_38[779]    = ( l_39 [779]);
assign l_38[780]    = ( l_39 [780]);
assign l_38[781]    = ( l_39 [781]);
assign l_38[782]    = ( l_39 [782]);
assign l_38[783]    = ( l_39 [783]);
assign l_38[784]    = ( l_39 [784]);
assign l_38[785]    = ( l_39 [785]);
assign l_38[786]    = ( l_39 [786]);
assign l_38[787]    = ( l_39 [787]);
assign l_38[788]    = ( l_39 [788]);
assign l_38[789]    = ( l_39 [789]);
assign l_38[790]    = ( l_39 [790]);
assign l_38[791]    = ( l_39 [791]);
assign l_38[792]    = ( l_39 [792]);
assign l_38[793]    = ( l_39 [793]);
assign l_38[794]    = ( l_39 [794]);
assign l_38[795]    = ( l_39 [795]);
assign l_38[796]    = ( l_39 [796]);
assign l_38[797]    = ( l_39 [797]);
assign l_38[798]    = ( l_39 [798]);
assign l_38[799]    = ( l_39 [799]);
assign l_38[800]    = ( l_39 [800]);
assign l_38[801]    = ( l_39 [801]);
assign l_38[802]    = ( l_39 [802]);
assign l_38[803]    = ( l_39 [803]);
assign l_38[804]    = ( l_39 [804]);
assign l_38[805]    = ( l_39 [805]);
assign l_38[806]    = ( l_39 [806]);
assign l_38[807]    = ( l_39 [807]);
assign l_38[808]    = ( l_39 [808]);
assign l_38[809]    = ( l_39 [809]);
assign l_38[810]    = ( l_39 [810]);
assign l_38[811]    = ( l_39 [811]);
assign l_38[812]    = ( l_39 [812]);
assign l_38[813]    = ( l_39 [813]);
assign l_38[814]    = ( l_39 [814]);
assign l_38[815]    = ( l_39 [815]);
assign l_38[816]    = ( l_39 [816]);
assign l_38[817]    = ( l_39 [817]);
assign l_38[818]    = ( l_39 [818]);
assign l_38[819]    = ( l_39 [819]);
assign l_38[820]    = ( l_39 [820]);
assign l_38[821]    = ( l_39 [821]);
assign l_38[822]    = ( l_39 [822]);
assign l_38[823]    = ( l_39 [823]);
assign l_38[824]    = ( l_39 [824]);
assign l_38[825]    = ( l_39 [825]);
assign l_38[826]    = ( l_39 [826]);
assign l_38[827]    = ( l_39 [827]);
assign l_38[828]    = ( l_39 [828]);
assign l_38[829]    = ( l_39 [829]);
assign l_38[830]    = ( l_39 [830]);
assign l_38[831]    = ( l_39 [831]);
assign l_38[832]    = ( l_39 [832]);
assign l_38[833]    = ( l_39 [833]);
assign l_38[834]    = ( l_39 [834]);
assign l_38[835]    = ( l_39 [835]);
assign l_38[836]    = ( l_39 [836]);
assign l_38[837]    = ( l_39 [837]);
assign l_38[838]    = ( l_39 [838]);
assign l_38[839]    = ( l_39 [839]);
assign l_38[840]    = ( l_39 [840]);
assign l_38[841]    = ( l_39 [841]);
assign l_38[842]    = ( l_39 [842]);
assign l_38[843]    = ( l_39 [843]);
assign l_38[844]    = ( l_39 [844]);
assign l_38[845]    = ( l_39 [845]);
assign l_38[846]    = ( l_39 [846]);
assign l_38[847]    = ( l_39 [847]);
assign l_38[848]    = ( l_39 [848]);
assign l_38[849]    = ( l_39 [849]);
assign l_38[850]    = ( l_39 [850]);
assign l_38[851]    = ( l_39 [851]);
assign l_38[852]    = ( l_39 [852]);
assign l_38[853]    = ( l_39 [853]);
assign l_38[854]    = ( l_39 [854]);
assign l_38[855]    = ( l_39 [855]);
assign l_38[856]    = ( l_39 [856]);
assign l_38[857]    = ( l_39 [857]);
assign l_38[858]    = ( l_39 [858]);
assign l_38[859]    = ( l_39 [859]);
assign l_38[860]    = ( l_39 [860]);
assign l_38[861]    = ( l_39 [861]);
assign l_38[862]    = ( l_39 [862]);
assign l_38[863]    = ( l_39 [863]);
assign l_38[864]    = ( l_39 [864]);
assign l_38[865]    = ( l_39 [865]);
assign l_38[866]    = ( l_39 [866]);
assign l_38[867]    = ( l_39 [867]);
assign l_38[868]    = ( l_39 [868]);
assign l_38[869]    = ( l_39 [869]);
assign l_38[870]    = ( l_39 [870]);
assign l_38[871]    = ( l_39 [871]);
assign l_38[872]    = ( l_39 [872]);
assign l_38[873]    = ( l_39 [873]);
assign l_38[874]    = ( l_39 [874]);
assign l_38[875]    = ( l_39 [875]);
assign l_38[876]    = ( l_39 [876]);
assign l_38[877]    = ( l_39 [877]);
assign l_38[878]    = ( l_39 [878]);
assign l_38[879]    = ( l_39 [879]);
assign l_38[880]    = ( l_39 [880]);
assign l_38[881]    = ( l_39 [881]);
assign l_38[882]    = ( l_39 [882]);
assign l_38[883]    = ( l_39 [883]);
assign l_38[884]    = ( l_39 [884]);
assign l_38[885]    = ( l_39 [885]);
assign l_38[886]    = ( l_39 [886]);
assign l_38[887]    = ( l_39 [887]);
assign l_38[888]    = ( l_39 [888]);
assign l_38[889]    = ( l_39 [889]);
assign l_38[890]    = ( l_39 [890]);
assign l_38[891]    = ( l_39 [891]);
assign l_38[892]    = ( l_39 [892]);
assign l_38[893]    = ( l_39 [893]);
assign l_38[894]    = ( l_39 [894]);
assign l_38[895]    = ( l_39 [895]);
assign l_38[896]    = ( l_39 [896]);
assign l_38[897]    = ( l_39 [897]);
assign l_38[898]    = ( l_39 [898]);
assign l_38[899]    = ( l_39 [899]);
assign l_38[900]    = ( l_39 [900]);
assign l_38[901]    = ( l_39 [901]);
assign l_38[902]    = ( l_39 [902]);
assign l_38[903]    = ( l_39 [903]);
assign l_38[904]    = ( l_39 [904]);
assign l_38[905]    = ( l_39 [905]);
assign l_38[906]    = ( l_39 [906]);
assign l_38[907]    = ( l_39 [907]);
assign l_38[908]    = ( l_39 [908]);
assign l_38[909]    = ( l_39 [909]);
assign l_38[910]    = ( l_39 [910]);
assign l_38[911]    = ( l_39 [911]);
assign l_38[912]    = ( l_39 [912]);
assign l_38[913]    = ( l_39 [913]);
assign l_38[914]    = ( l_39 [914]);
assign l_38[915]    = ( l_39 [915]);
assign l_38[916]    = ( l_39 [916]);
assign l_38[917]    = ( l_39 [917]);
assign l_38[918]    = ( l_39 [918]);
assign l_38[919]    = ( l_39 [919]);
assign l_38[920]    = ( l_39 [920]);
assign l_38[921]    = ( l_39 [921]);
assign l_38[922]    = ( l_39 [922]);
assign l_38[923]    = ( l_39 [923]);
assign l_38[924]    = ( l_39 [924]);
assign l_38[925]    = ( l_39 [925]);
assign l_38[926]    = ( l_39 [926]);
assign l_38[927]    = ( l_39 [927]);
assign l_38[928]    = ( l_39 [928]);
assign l_38[929]    = ( l_39 [929]);
assign l_38[930]    = ( l_39 [930]);
assign l_38[931]    = ( l_39 [931]);
assign l_38[932]    = ( l_39 [932]);
assign l_38[933]    = ( l_39 [933]);
assign l_38[934]    = ( l_39 [934]);
assign l_38[935]    = ( l_39 [935]);
assign l_38[936]    = ( l_39 [936]);
assign l_38[937]    = ( l_39 [937]);
assign l_38[938]    = ( l_39 [938]);
assign l_38[939]    = ( l_39 [939]);
assign l_38[940]    = ( l_39 [940]);
assign l_38[941]    = ( l_39 [941]);
assign l_38[942]    = ( l_39 [942]);
assign l_38[943]    = ( l_39 [943]);
assign l_38[944]    = ( l_39 [944]);
assign l_38[945]    = ( l_39 [945]);
assign l_38[946]    = ( l_39 [946]);
assign l_38[947]    = ( l_39 [947]);
assign l_38[948]    = ( l_39 [948]);
assign l_38[949]    = ( l_39 [949]);
assign l_38[950]    = ( l_39 [950]);
assign l_38[951]    = ( l_39 [951]);
assign l_38[952]    = ( l_39 [952]);
assign l_38[953]    = ( l_39 [953]);
assign l_38[954]    = ( l_39 [954]);
assign l_38[955]    = ( l_39 [955]);
assign l_38[956]    = ( l_39 [956]);
assign l_38[957]    = ( l_39 [957]);
assign l_38[958]    = ( l_39 [958]);
assign l_38[959]    = ( l_39 [959]);
assign l_38[960]    = ( l_39 [960]);
assign l_38[961]    = ( l_39 [961]);
assign l_38[962]    = ( l_39 [962]);
assign l_38[963]    = ( l_39 [963]);
assign l_38[964]    = ( l_39 [964]);
assign l_38[965]    = ( l_39 [965]);
assign l_38[966]    = ( l_39 [966]);
assign l_38[967]    = ( l_39 [967]);
assign l_38[968]    = ( l_39 [968]);
assign l_38[969]    = ( l_39 [969]);
assign l_38[970]    = ( l_39 [970]);
assign l_38[971]    = ( l_39 [971]);
assign l_38[972]    = ( l_39 [972]);
assign l_38[973]    = ( l_39 [973]);
assign l_38[974]    = ( l_39 [974]);
assign l_38[975]    = ( l_39 [975]);
assign l_38[976]    = ( l_39 [976]);
assign l_38[977]    = ( l_39 [977]);
assign l_38[978]    = ( l_39 [978]);
assign l_38[979]    = ( l_39 [979]);
assign l_38[980]    = ( l_39 [980]);
assign l_38[981]    = ( l_39 [981]);
assign l_38[982]    = ( l_39 [982]);
assign l_38[983]    = ( l_39 [983]);
assign l_38[984]    = ( l_39 [984]);
assign l_38[985]    = ( l_39 [985]);
assign l_38[986]    = ( l_39 [986]);
assign l_38[987]    = ( l_39 [987]);
assign l_38[988]    = ( l_39 [988]);
assign l_38[989]    = ( l_39 [989]);
assign l_38[990]    = ( l_39 [990]);
assign l_38[991]    = ( l_39 [991]);
assign l_38[992]    = ( l_39 [992]);
assign l_38[993]    = ( l_39 [993]);
assign l_38[994]    = ( l_39 [994]);
assign l_38[995]    = ( l_39 [995]);
assign l_38[996]    = ( l_39 [996]);
assign l_38[997]    = ( l_39 [997]);
assign l_38[998]    = ( l_39 [998]);
assign l_38[999]    = ( l_39 [999]);
assign l_38[1000]    = ( l_39 [1000]);
assign l_38[1001]    = ( l_39 [1001]);
assign l_38[1002]    = ( l_39 [1002]);
assign l_38[1003]    = ( l_39 [1003]);
assign l_38[1004]    = ( l_39 [1004]);
assign l_38[1005]    = ( l_39 [1005]);
assign l_38[1006]    = ( l_39 [1006]);
assign l_38[1007]    = ( l_39 [1007]);
assign l_38[1008]    = ( l_39 [1008]);
assign l_38[1009]    = ( l_39 [1009]);
assign l_38[1010]    = ( l_39 [1010]);
assign l_38[1011]    = ( l_39 [1011]);
assign l_38[1012]    = ( l_39 [1012]);
assign l_38[1013]    = ( l_39 [1013]);
assign l_38[1014]    = ( l_39 [1014]);
assign l_38[1015]    = ( l_39 [1015]);
assign l_38[1016]    = ( l_39 [1016]);
assign l_38[1017]    = ( l_39 [1017]);
assign l_38[1018]    = ( l_39 [1018]);
assign l_38[1019]    = ( l_39 [1019]);
assign l_38[1020]    = ( l_39 [1020]);
assign l_38[1021]    = ( l_39 [1021]);
assign l_38[1022]    = ( l_39 [1022]);
assign l_38[1023]    = ( l_39 [1023]);
assign l_38[1024]    = ( l_39 [1024]);
assign l_38[1025]    = ( l_39 [1025]);
assign l_38[1026]    = ( l_39 [1026]);
assign l_38[1027]    = ( l_39 [1027]);
assign l_38[1028]    = ( l_39 [1028]);
assign l_38[1029]    = ( l_39 [1029]);
assign l_38[1030]    = ( l_39 [1030]);
assign l_38[1031]    = ( l_39 [1031]);
assign l_38[1032]    = ( l_39 [1032]);
assign l_38[1033]    = ( l_39 [1033]);
assign l_38[1034]    = ( l_39 [1034]);
assign l_38[1035]    = ( l_39 [1035]);
assign l_38[1036]    = ( l_39 [1036]);
assign l_38[1037]    = ( l_39 [1037]);
assign l_38[1038]    = ( l_39 [1038]);
assign l_38[1039]    = ( l_39 [1039]);
assign l_38[1040]    = ( l_39 [1040]);
assign l_38[1041]    = ( l_39 [1041]);
assign l_38[1042]    = ( l_39 [1042] & !i[1814]) | ( l_39 [1043] &  i[1814]);
assign l_38[1043]    = ( l_39 [1044] & !i[1814]) | ( l_39 [1045] &  i[1814]);
assign l_38[1044]    = ( l_39 [1046] & !i[1814]) | ( l_39 [1047] &  i[1814]);
assign l_38[1045]    = ( l_39 [1048] & !i[1814]) | ( l_39 [1049] &  i[1814]);
assign l_38[1046]    = ( l_39 [1050] & !i[1814]) | ( l_39 [1051] &  i[1814]);
assign l_38[1047]    = ( l_39 [1052] & !i[1814]) | ( l_39 [1053] &  i[1814]);
assign l_38[1048]    = ( l_39 [1054] & !i[1814]) | ( l_39 [1055] &  i[1814]);
assign l_38[1049]    = ( l_39 [1056] & !i[1814]) | ( l_39 [1057] &  i[1814]);
assign l_38[1050]    = ( l_39 [1058] & !i[1814]) | ( l_39 [1059] &  i[1814]);
assign l_38[1051]    = ( l_39 [1060] & !i[1814]) | ( l_39 [1061] &  i[1814]);
assign l_38[1052]    = ( l_39 [1062] & !i[1814]) | ( l_39 [1063] &  i[1814]);
assign l_38[1053]    = ( l_39 [1064] & !i[1814]) | ( l_39 [1065] &  i[1814]);
assign l_38[1054]    = ( l_39 [1066] & !i[1814]) | ( l_39 [1067] &  i[1814]);
assign l_38[1055]    = ( l_39 [1068] & !i[1814]) | ( l_39 [1069] &  i[1814]);
assign l_38[1056]    = ( l_39 [1070] & !i[1814]) | ( l_39 [1071] &  i[1814]);
assign l_38[1057]    = ( l_39 [1072] & !i[1814]) | ( l_39 [1073] &  i[1814]);
assign l_38[1058]    = ( l_39 [1074] & !i[1814]) | ( l_39 [1075] &  i[1814]);
assign l_38[1059]    = ( l_39 [1076] & !i[1814]) | ( l_39 [1077] &  i[1814]);
assign l_38[1060]    = ( l_39 [1078] & !i[1814]) | ( l_39 [1079] &  i[1814]);
assign l_38[1061]    = ( l_39 [1080] & !i[1814]) | ( l_39 [1081] &  i[1814]);
assign l_38[1062]    = ( l_39 [1082] & !i[1814]) | ( l_39 [1083] &  i[1814]);
assign l_38[1063]    = ( l_39 [1084] & !i[1814]) | ( l_39 [1085] &  i[1814]);
assign l_38[1064]    = ( l_39 [1086] & !i[1814]) | ( l_39 [1087] &  i[1814]);
assign l_38[1065]    = ( l_39 [1088] & !i[1814]) | ( l_39 [1089] &  i[1814]);
assign l_38[1066]    = ( l_39 [1090] & !i[1814]) | ( l_39 [1091] &  i[1814]);
assign l_38[1067]    = ( l_39 [1092] & !i[1814]) | ( l_39 [1093] &  i[1814]);
assign l_38[1068]    = ( l_39 [1094] & !i[1814]) | ( l_39 [1095] &  i[1814]);
assign l_38[1069]    = ( l_39 [1096] & !i[1814]) | ( l_39 [1097] &  i[1814]);
assign l_38[1070]    = ( l_39 [1098] & !i[1814]) | ( l_39 [1099] &  i[1814]);
assign l_38[1071]    = ( l_39 [1100] & !i[1814]) | ( l_39 [1101] &  i[1814]);
assign l_38[1072]    = ( l_39 [1102] & !i[1814]) | ( l_39 [1103] &  i[1814]);
assign l_38[1073]    = ( l_39 [1104] & !i[1814]) | ( l_39 [1105] &  i[1814]);
assign l_38[1074]    = ( l_39 [1106] & !i[1814]) | ( l_39 [1107] &  i[1814]);
assign l_38[1075]    = ( l_39 [1108] & !i[1814]) | ( l_39 [1109] &  i[1814]);
assign l_38[1076]    = ( l_39 [1110] & !i[1814]) | ( l_39 [1111] &  i[1814]);
assign l_38[1077]    = ( l_39 [1112] & !i[1814]) | ( l_39 [1113] &  i[1814]);
assign l_38[1078]    = ( l_39 [1114] & !i[1814]) | ( l_39 [1115] &  i[1814]);
assign l_38[1079]    = ( l_39 [1116] & !i[1814]) | ( l_39 [1117] &  i[1814]);
assign l_38[1080]    = ( l_39 [1118] & !i[1814]) | ( l_39 [1119] &  i[1814]);
assign l_38[1081]    = ( l_39 [1120] & !i[1814]) | ( l_39 [1121] &  i[1814]);
assign l_38[1082]    = ( l_39 [1122] & !i[1814]) | ( l_39 [1123] &  i[1814]);
assign l_38[1083]    = ( l_39 [1124] & !i[1814]) | ( l_39 [1125] &  i[1814]);
assign l_38[1084]    = ( l_39 [1126] & !i[1814]) | ( l_39 [1127] &  i[1814]);
assign l_38[1085]    = ( l_39 [1128] & !i[1814]) | ( l_39 [1129] &  i[1814]);
assign l_38[1086]    = ( l_39 [1130] & !i[1814]) | ( l_39 [1131] &  i[1814]);
assign l_38[1087]    = ( l_39 [1132] & !i[1814]) | ( l_39 [1133] &  i[1814]);
assign l_38[1088]    = ( l_39 [1134] & !i[1814]) | ( l_39 [1135] &  i[1814]);
assign l_38[1089]    = ( l_39 [1136] & !i[1814]) | ( l_39 [1137] &  i[1814]);
assign l_38[1090]    = ( l_39 [1138] & !i[1814]) | ( l_39 [1139] &  i[1814]);
assign l_38[1091]    = ( l_39 [1140] & !i[1814]) | ( l_39 [1141] &  i[1814]);
assign l_38[1092]    = ( l_39 [1142] & !i[1814]) | ( l_39 [1143] &  i[1814]);
assign l_38[1093]    = ( l_39 [1144] & !i[1814]) | ( l_39 [1145] &  i[1814]);
assign l_38[1094]    = ( l_39 [1146] & !i[1814]) | ( l_39 [1147] &  i[1814]);
assign l_38[1095]    = ( l_39 [1148] & !i[1814]) | ( l_39 [1149] &  i[1814]);
assign l_38[1096]    = ( l_39 [1150] & !i[1814]) | ( l_39 [1151] &  i[1814]);
assign l_38[1097]    = ( l_39 [1152] & !i[1814]) | ( l_39 [1153] &  i[1814]);
assign l_38[1098]    = ( l_39 [1154] & !i[1814]) | ( l_39 [1155] &  i[1814]);
assign l_38[1099]    = ( l_39 [1156] & !i[1814]) | ( l_39 [1157] &  i[1814]);
assign l_38[1100]    = ( l_39 [1158] & !i[1814]) | ( l_39 [1159] &  i[1814]);
assign l_38[1101]    = ( l_39 [1160] & !i[1814]) | ( l_39 [1161] &  i[1814]);
assign l_38[1102]    = ( l_39 [1162] & !i[1814]) | ( l_39 [1163] &  i[1814]);
assign l_38[1103]    = ( l_39 [1164] & !i[1814]) | ( l_39 [1165] &  i[1814]);
assign l_38[1104]    = ( l_39 [1166] & !i[1814]) | ( l_39 [1167] &  i[1814]);
assign l_38[1105]    = ( l_39 [1168] & !i[1814]) | ( l_39 [1169] &  i[1814]);
assign l_38[1106]    = ( l_39 [1170] & !i[1814]) | ( l_39 [1171] &  i[1814]);
assign l_38[1107]    = ( l_39 [1172] & !i[1814]) | ( l_39 [1173] &  i[1814]);
assign l_38[1108]    = ( l_39 [1174] & !i[1814]) | ( l_39 [1175] &  i[1814]);
assign l_38[1109]    = ( l_39 [1176] & !i[1814]) | ( l_39 [1177] &  i[1814]);
assign l_38[1110]    = ( l_39 [1178] & !i[1814]) | ( l_39 [1179] &  i[1814]);
assign l_38[1111]    = ( l_39 [1180] & !i[1814]) | ( l_39 [1181] &  i[1814]);
assign l_38[1112]    = ( l_39 [1182] & !i[1814]) | ( l_39 [1183] &  i[1814]);
assign l_38[1113]    = ( l_39 [1184] & !i[1814]) | ( l_39 [1185] &  i[1814]);
assign l_38[1114]    = ( l_39 [1186] & !i[1814]) | ( l_39 [1187] &  i[1814]);
assign l_38[1115]    = ( l_39 [1188] & !i[1814]) | ( l_39 [1189] &  i[1814]);
assign l_38[1116]    = ( l_39 [1190] & !i[1814]) | ( l_39 [1191] &  i[1814]);
assign l_38[1117]    = ( l_39 [1192] & !i[1814]) | ( l_39 [1193] &  i[1814]);
assign l_38[1118]    = ( l_39 [1194] & !i[1814]) | ( l_39 [1195] &  i[1814]);
assign l_38[1119]    = ( l_39 [1196] & !i[1814]) | ( l_39 [1197] &  i[1814]);
assign l_38[1120]    = ( l_39 [1198] & !i[1814]) | ( l_39 [1199] &  i[1814]);
assign l_38[1121]    = ( l_39 [1200] & !i[1814]) | ( l_39 [1201] &  i[1814]);
assign l_38[1122]    = ( l_39 [1202] & !i[1814]) | ( l_39 [1203] &  i[1814]);
assign l_38[1123]    = ( l_39 [1204] & !i[1814]) | ( l_39 [1205] &  i[1814]);
assign l_38[1124]    = ( l_39 [1206] & !i[1814]) | ( l_39 [1207] &  i[1814]);
assign l_38[1125]    = ( l_39 [1208] & !i[1814]) | ( l_39 [1209] &  i[1814]);
assign l_38[1126]    = ( l_39 [1210] & !i[1814]) | ( l_39 [1211] &  i[1814]);
assign l_38[1127]    = ( l_39 [1212] & !i[1814]) | ( l_39 [1213] &  i[1814]);
assign l_38[1128]    = ( l_39 [1214] & !i[1814]) | ( l_39 [1215] &  i[1814]);
assign l_38[1129]    = ( l_39 [1216] & !i[1814]) | ( l_39 [1217] &  i[1814]);
assign l_38[1130]    = ( l_39 [1218] & !i[1814]) | ( l_39 [1219] &  i[1814]);
assign l_38[1131]    = ( l_39 [1220] & !i[1814]) | ( l_39 [1221] &  i[1814]);
assign l_38[1132]    = ( l_39 [1222] & !i[1814]) | ( l_39 [1223] &  i[1814]);
assign l_38[1133]    = ( l_39 [1224] & !i[1814]) | ( l_39 [1225] &  i[1814]);
assign l_38[1134]    = ( l_39 [1226] & !i[1814]) | ( l_39 [1227] &  i[1814]);
assign l_38[1135]    = ( l_39 [1228] & !i[1814]) | ( l_39 [1229] &  i[1814]);
assign l_38[1136]    = ( l_39 [1230] & !i[1814]) | ( l_39 [1231] &  i[1814]);
assign l_38[1137]    = ( l_39 [1232] & !i[1814]) | ( l_39 [1233] &  i[1814]);
assign l_38[1138]    = ( l_39 [1234] & !i[1814]) | ( l_39 [1235] &  i[1814]);
assign l_38[1139]    = ( l_39 [1236] & !i[1814]) | ( l_39 [1237] &  i[1814]);
assign l_38[1140]    = ( l_39 [1238] & !i[1814]) | ( l_39 [1239] &  i[1814]);
assign l_38[1141]    = ( l_39 [1240] & !i[1814]) | ( l_39 [1241] &  i[1814]);
assign l_38[1142]    = ( l_39 [1242] & !i[1814]) | ( l_39 [1243] &  i[1814]);
assign l_38[1143]    = ( l_39 [1244] & !i[1814]) | ( l_39 [1245] &  i[1814]);
assign l_38[1144]    = ( l_39 [1246] & !i[1814]) | ( l_39 [1247] &  i[1814]);
assign l_38[1145]    = ( l_39 [1248] & !i[1814]) | ( l_39 [1249] &  i[1814]);
assign l_38[1146]    = ( l_39 [1250] & !i[1814]) | ( l_39 [1251] &  i[1814]);
assign l_38[1147]    = ( l_39 [1252] & !i[1814]) | ( l_39 [1253] &  i[1814]);
assign l_38[1148]    = ( l_39 [1254] & !i[1814]) | ( l_39 [1255] &  i[1814]);
assign l_38[1149]    = ( l_39 [1256] & !i[1814]) | ( l_39 [1257] &  i[1814]);
assign l_38[1150]    = ( l_39 [1258] & !i[1814]) | ( l_39 [1259] &  i[1814]);
assign l_38[1151]    = ( l_39 [1260] & !i[1814]) | ( l_39 [1261] &  i[1814]);
assign l_38[1152]    = ( l_39 [1262] & !i[1814]) | ( l_39 [1263] &  i[1814]);
assign l_38[1153]    = ( l_39 [1264] & !i[1814]) | ( l_39 [1265] &  i[1814]);
assign l_38[1154]    = ( l_39 [1266] & !i[1814]) | ( l_39 [1267] &  i[1814]);
assign l_38[1155]    = ( l_39 [1268] & !i[1814]) | ( l_39 [1269] &  i[1814]);
assign l_38[1156]    = ( l_39 [1270] & !i[1814]) | ( l_39 [1271] &  i[1814]);
assign l_38[1157]    = ( l_39 [1272] & !i[1814]) | ( l_39 [1273] &  i[1814]);
assign l_38[1158]    = ( l_39 [1274] & !i[1814]) | ( l_39 [1275] &  i[1814]);
assign l_38[1159]    = ( l_39 [1276] & !i[1814]) | ( l_39 [1277] &  i[1814]);
assign l_38[1160]    = ( l_39 [1278] & !i[1814]) | ( l_39 [1279] &  i[1814]);
assign l_38[1161]    = ( l_39 [1280] & !i[1814]) | ( l_39 [1281] &  i[1814]);
assign l_38[1162]    = ( l_39 [1282] & !i[1814]) | ( l_39 [1283] &  i[1814]);
assign l_38[1163]    = ( l_39 [1284] & !i[1814]) | ( l_39 [1285] &  i[1814]);
assign l_38[1164]    = ( l_39 [1286] & !i[1814]) | ( l_39 [1287] &  i[1814]);
assign l_38[1165]    = ( l_39 [1288] & !i[1814]) | ( l_39 [1289] &  i[1814]);
assign l_38[1166]    = ( l_39 [1290] & !i[1814]) | ( l_39 [1291] &  i[1814]);
assign l_38[1167]    = ( l_39 [1292] & !i[1814]) | ( l_39 [1293] &  i[1814]);
assign l_38[1168]    = ( l_39 [1294] & !i[1814]) | ( l_39 [1295] &  i[1814]);
assign l_38[1169]    = ( l_39 [1296] & !i[1814]) | ( l_39 [1297] &  i[1814]);
assign l_38[1170]    = ( l_39 [1298] & !i[1814]) | ( l_39 [1299] &  i[1814]);
assign l_38[1171]    = ( l_39 [1300] & !i[1814]) | ( l_39 [1301] &  i[1814]);
assign l_38[1172]    = ( l_39 [1302] & !i[1814]) | ( l_39 [1303] &  i[1814]);
assign l_38[1173]    = ( l_39 [1304] & !i[1814]) | ( l_39 [1305] &  i[1814]);
assign l_38[1174]    = ( l_39 [1306] & !i[1814]) | ( l_39 [1307] &  i[1814]);
assign l_38[1175]    = ( l_39 [1308] & !i[1814]) | ( l_39 [1309] &  i[1814]);
assign l_38[1176]    = ( l_39 [1310] & !i[1814]) | ( l_39 [1311] &  i[1814]);
assign l_38[1177]    = ( l_39 [1312] & !i[1814]) | ( l_39 [1313] &  i[1814]);
assign l_38[1178]    = ( l_39 [1314] & !i[1814]) | ( l_39 [1315] &  i[1814]);
assign l_38[1179]    = ( l_39 [1316] & !i[1814]) | ( l_39 [1317] &  i[1814]);
assign l_38[1180]    = ( l_39 [1318] & !i[1814]) | ( l_39 [1319] &  i[1814]);
assign l_38[1181]    = ( l_39 [1320] & !i[1814]) | ( l_39 [1321] &  i[1814]);
assign l_38[1182]    = ( l_39 [1322] & !i[1814]) | ( l_39 [1323] &  i[1814]);
assign l_38[1183]    = ( l_39 [1324] & !i[1814]) | ( l_39 [1325] &  i[1814]);
assign l_38[1184]    = ( l_39 [1326] & !i[1814]) | ( l_39 [1327] &  i[1814]);
assign l_38[1185]    = ( l_39 [1328] & !i[1814]) | ( l_39 [1329] &  i[1814]);
assign l_38[1186]    = ( l_39 [1330] & !i[1814]) | ( l_39 [1331] &  i[1814]);
assign l_38[1187]    = ( l_39 [1332] & !i[1814]) | ( l_39 [1333] &  i[1814]);
assign l_38[1188]    = ( l_39 [1334] & !i[1814]) | ( l_39 [1335] &  i[1814]);
assign l_38[1189]    = ( l_39 [1336] & !i[1814]) | ( l_39 [1337] &  i[1814]);
assign l_38[1190]    = ( l_39 [1338] & !i[1814]) | ( l_39 [1339] &  i[1814]);
assign l_38[1191]    = ( l_39 [1340] & !i[1814]) | ( l_39 [1341] &  i[1814]);
assign l_38[1192]    = ( l_39 [1342] & !i[1814]) | ( l_39 [1343] &  i[1814]);
assign l_38[1193]    = ( l_39 [1344] & !i[1814]) | ( l_39 [1345] &  i[1814]);
assign l_38[1194]    = ( l_39 [1346] & !i[1814]) | ( l_39 [1347] &  i[1814]);
assign l_38[1195]    = ( l_39 [1348] & !i[1814]) | ( l_39 [1349] &  i[1814]);
assign l_38[1196]    = ( l_39 [1350] & !i[1814]) | ( l_39 [1351] &  i[1814]);
assign l_38[1197]    = ( l_39 [1352] & !i[1814]) | ( l_39 [1353] &  i[1814]);
assign l_38[1198]    = ( l_39 [1354] & !i[1814]) | ( l_39 [1355] &  i[1814]);
assign l_38[1199]    = ( l_39 [1356] & !i[1814]) | ( l_39 [1357] &  i[1814]);
assign l_38[1200]    = ( l_39 [1358] & !i[1814]) | ( l_39 [1359] &  i[1814]);
assign l_38[1201]    = ( l_39 [1360] & !i[1814]) | ( l_39 [1361] &  i[1814]);
assign l_38[1202]    = ( l_39 [1362] & !i[1814]) | ( l_39 [1363] &  i[1814]);
assign l_38[1203]    = ( l_39 [1364] & !i[1814]) | ( l_39 [1365] &  i[1814]);
assign l_38[1204]    = ( l_39 [1366] & !i[1814]) | ( l_39 [1367] &  i[1814]);
assign l_38[1205]    = ( l_39 [1368] & !i[1814]) | ( l_39 [1369] &  i[1814]);
assign l_38[1206]    = ( l_39 [1370] & !i[1814]) | ( l_39 [1371] &  i[1814]);
assign l_38[1207]    = ( l_39 [1372] & !i[1814]) | ( l_39 [1373] &  i[1814]);
assign l_38[1208]    = ( l_39 [1374] & !i[1814]) | ( l_39 [1375] &  i[1814]);
assign l_38[1209]    = ( l_39 [1376] & !i[1814]) | ( l_39 [1377] &  i[1814]);
assign l_38[1210]    = ( l_39 [1378] & !i[1814]) | ( l_39 [1379] &  i[1814]);
assign l_38[1211]    = ( l_39 [1380] & !i[1814]) | ( l_39 [1381] &  i[1814]);
assign l_38[1212]    = ( l_39 [1382] & !i[1814]) | ( l_39 [1383] &  i[1814]);
assign l_38[1213]    = ( l_39 [1384] & !i[1814]) | ( l_39 [1385] &  i[1814]);
assign l_38[1214]    = ( l_39 [1386] & !i[1814]) | ( l_39 [1387] &  i[1814]);
assign l_38[1215]    = ( l_39 [1388] & !i[1814]) | ( l_39 [1389] &  i[1814]);
assign l_38[1216]    = ( l_39 [1390] & !i[1814]) | ( l_39 [1391] &  i[1814]);
assign l_38[1217]    = ( l_39 [1392] & !i[1814]) | ( l_39 [1393] &  i[1814]);
assign l_38[1218]    = ( l_39 [1394] & !i[1814]) | ( l_39 [1395] &  i[1814]);
assign l_38[1219]    = ( l_39 [1396] & !i[1814]) | ( l_39 [1397] &  i[1814]);
assign l_38[1220]    = ( l_39 [1398] & !i[1814]) | ( l_39 [1399] &  i[1814]);
assign l_38[1221]    = ( l_39 [1400] & !i[1814]) | ( l_39 [1401] &  i[1814]);
assign l_38[1222]    = ( l_39 [1402] & !i[1814]) | ( l_39 [1403] &  i[1814]);
assign l_38[1223]    = ( l_39 [1404] & !i[1814]) | ( l_39 [1405] &  i[1814]);
assign l_38[1224]    = ( l_39 [1406] & !i[1814]) | ( l_39 [1407] &  i[1814]);
assign l_38[1225]    = ( l_39 [1408] & !i[1814]) | ( l_39 [1409] &  i[1814]);
assign l_38[1226]    = ( l_39 [1410] & !i[1814]) | ( l_39 [1411] &  i[1814]);
assign l_38[1227]    = ( l_39 [1412] & !i[1814]) | ( l_39 [1413] &  i[1814]);
assign l_38[1228]    = ( l_39 [1414] & !i[1814]) | ( l_39 [1415] &  i[1814]);
assign l_38[1229]    = ( l_39 [1416] & !i[1814]) | ( l_39 [1417] &  i[1814]);
assign l_38[1230]    = ( l_39 [1418] & !i[1814]) | ( l_39 [1419] &  i[1814]);
assign l_38[1231]    = ( l_39 [1420] & !i[1814]) | ( l_39 [1421] &  i[1814]);
assign l_38[1232]    = ( l_39 [1422] & !i[1814]) | ( l_39 [1423] &  i[1814]);
assign l_38[1233]    = ( l_39 [1424] & !i[1814]) | ( l_39 [1425] &  i[1814]);
assign l_38[1234]    = ( l_39 [1426] & !i[1814]) | ( l_39 [1427] &  i[1814]);
assign l_38[1235]    = ( l_39 [1428] & !i[1814]) | ( l_39 [1429] &  i[1814]);
assign l_38[1236]    = ( l_39 [1430] & !i[1814]) | ( l_39 [1431] &  i[1814]);
assign l_38[1237]    = ( l_39 [1432] & !i[1814]) | ( l_39 [1433] &  i[1814]);
assign l_38[1238]    = ( l_39 [1434] & !i[1814]) | ( l_39 [1435] &  i[1814]);
assign l_38[1239]    = ( l_39 [1436] & !i[1814]) | ( l_39 [1437] &  i[1814]);
assign l_38[1240]    = ( l_39 [1438] & !i[1814]) | ( l_39 [1439] &  i[1814]);
assign l_38[1241]    = ( l_39 [1440] & !i[1814]) | ( l_39 [1441] &  i[1814]);
assign l_38[1242]    = ( l_39 [1442] & !i[1814]) | ( l_39 [1443] &  i[1814]);
assign l_38[1243]    = ( l_39 [1444] & !i[1814]) | ( l_39 [1445] &  i[1814]);
assign l_38[1244]    = ( l_39 [1446] & !i[1814]) | ( l_39 [1447] &  i[1814]);
assign l_38[1245]    = ( l_39 [1448] & !i[1814]) | ( l_39 [1449] &  i[1814]);
assign l_38[1246]    = ( l_39 [1450] & !i[1814]) | ( l_39 [1451] &  i[1814]);
assign l_38[1247]    = ( l_39 [1452] & !i[1814]) | ( l_39 [1453] &  i[1814]);
assign l_38[1248]    = ( l_39 [1454] & !i[1814]) | ( l_39 [1455] &  i[1814]);
assign l_38[1249]    = ( l_39 [1456] & !i[1814]) | ( l_39 [1457] &  i[1814]);
assign l_38[1250]    = ( l_39 [1458] & !i[1814]) | ( l_39 [1459] &  i[1814]);
assign l_38[1251]    = ( l_39 [1460] & !i[1814]) | ( l_39 [1461] &  i[1814]);
assign l_38[1252]    = ( l_39 [1462] & !i[1814]) | ( l_39 [1463] &  i[1814]);
assign l_38[1253]    = ( l_39 [1464] & !i[1814]) | ( l_39 [1465] &  i[1814]);
assign l_38[1254]    = ( l_39 [1466] & !i[1814]) | ( l_39 [1467] &  i[1814]);
assign l_38[1255]    = ( l_39 [1468] & !i[1814]) | ( l_39 [1469] &  i[1814]);
assign l_38[1256]    = ( l_39 [1470] & !i[1814]) | ( l_39 [1471] &  i[1814]);
assign l_38[1257]    = ( l_39 [1472] & !i[1814]) | ( l_39 [1473] &  i[1814]);
assign l_38[1258]    = ( l_39 [1474] & !i[1814]) | ( l_39 [1475] &  i[1814]);
assign l_38[1259]    = ( l_39 [1476] & !i[1814]) | ( l_39 [1477] &  i[1814]);
assign l_38[1260]    = ( l_39 [1478] & !i[1814]) | ( l_39 [1479] &  i[1814]);
assign l_38[1261]    = ( l_39 [1480] & !i[1814]) | ( l_39 [1481] &  i[1814]);
assign l_38[1262]    = ( l_39 [1482] & !i[1814]) | ( l_39 [1483] &  i[1814]);
assign l_38[1263]    = ( l_39 [1484] & !i[1814]) | ( l_39 [1485] &  i[1814]);
assign l_38[1264]    = ( l_39 [1486] & !i[1814]) | ( l_39 [1487] &  i[1814]);
assign l_38[1265]    = ( l_39 [1488] & !i[1814]) | ( l_39 [1489] &  i[1814]);
assign l_38[1266]    = ( l_39 [1490] & !i[1814]) | ( l_39 [1491] &  i[1814]);
assign l_38[1267]    = ( l_39 [1492] & !i[1814]) | ( l_39 [1493] &  i[1814]);
assign l_38[1268]    = ( l_39 [1494] & !i[1814]) | ( l_39 [1495] &  i[1814]);
assign l_38[1269]    = ( l_39 [1496] & !i[1814]) | ( l_39 [1497] &  i[1814]);
assign l_38[1270]    = ( l_39 [1498] & !i[1814]) | ( l_39 [1499] &  i[1814]);
assign l_38[1271]    = ( l_39 [1500] & !i[1814]) | ( l_39 [1501] &  i[1814]);
assign l_38[1272]    = ( l_39 [1502] & !i[1814]) | ( l_39 [1503] &  i[1814]);
assign l_38[1273]    = ( l_39 [1504] & !i[1814]) | ( l_39 [1505] &  i[1814]);
assign l_38[1274]    = ( l_39 [1506] & !i[1814]) | ( l_39 [1507] &  i[1814]);
assign l_38[1275]    = ( l_39 [1508] & !i[1814]) | ( l_39 [1509] &  i[1814]);
assign l_38[1276]    = ( l_39 [1510] & !i[1814]) | ( l_39 [1511] &  i[1814]);
assign l_38[1277]    = ( l_39 [1512] & !i[1814]) | ( l_39 [1513] &  i[1814]);
assign l_38[1278]    = ( l_39 [1514] & !i[1814]) | ( l_39 [1515] &  i[1814]);
assign l_38[1279]    = ( l_39 [1516] & !i[1814]) | ( l_39 [1517] &  i[1814]);
assign l_38[1280]    = ( l_39 [1518] & !i[1814]) | ( l_39 [1519] &  i[1814]);
assign l_38[1281]    = ( l_39 [1520] & !i[1814]) | ( l_39 [1521] &  i[1814]);
assign l_38[1282]    = ( l_39 [1522] & !i[1814]) | ( l_39 [1523] &  i[1814]);
assign l_38[1283]    = ( l_39 [1524] & !i[1814]) | ( l_39 [1525] &  i[1814]);
assign l_38[1284]    = ( l_39 [1526] & !i[1814]) | ( l_39 [1527] &  i[1814]);
assign l_38[1285]    = ( l_39 [1528] & !i[1814]) | ( l_39 [1529] &  i[1814]);
assign l_38[1286]    = ( l_39 [1530] & !i[1814]) | ( l_39 [1531] &  i[1814]);
assign l_38[1287]    = ( l_39 [1532] & !i[1814]) | ( l_39 [1533] &  i[1814]);
assign l_38[1288]    = ( l_39 [1534] & !i[1814]) | ( l_39 [1535] &  i[1814]);
assign l_38[1289]    = ( l_39 [1536] & !i[1814]) | ( l_39 [1537] &  i[1814]);
assign l_38[1290]    = ( l_39 [1538] & !i[1814]) | ( l_39 [1539] &  i[1814]);
assign l_38[1291]    = ( l_39 [1540] & !i[1814]) | ( l_39 [1541] &  i[1814]);
assign l_38[1292]    = ( l_39 [1542] & !i[1814]) | ( l_39 [1543] &  i[1814]);
assign l_38[1293]    = ( l_39 [1544] & !i[1814]) | ( l_39 [1545] &  i[1814]);
assign l_38[1294]    = ( l_39 [1546] & !i[1814]) | ( l_39 [1547] &  i[1814]);
assign l_38[1295]    = ( l_39 [1548] & !i[1814]) | ( l_39 [1549] &  i[1814]);
assign l_38[1296]    = ( l_39 [1550] & !i[1814]) | ( l_39 [1551] &  i[1814]);
assign l_38[1297]    = ( l_39 [1552] & !i[1814]) | ( l_39 [1553] &  i[1814]);
assign l_38[1298]    = ( l_39 [1554] & !i[1814]) | ( l_39 [1555] &  i[1814]);
assign l_38[1299]    = ( l_39 [1556] & !i[1814]) | ( l_39 [1557] &  i[1814]);
assign l_38[1300]    = ( l_39 [1558] & !i[1814]) | ( l_39 [1559] &  i[1814]);
assign l_38[1301]    = ( l_39 [1560] & !i[1814]) | ( l_39 [1561] &  i[1814]);
assign l_38[1302]    = ( l_39 [1562] & !i[1814]) | ( l_39 [1563] &  i[1814]);
assign l_38[1303]    = ( l_39 [1564] & !i[1814]) | ( l_39 [1565] &  i[1814]);
assign l_38[1304]    = ( l_39 [1566] & !i[1814]) | ( l_39 [1567] &  i[1814]);
assign l_38[1305]    = ( l_39 [1568] & !i[1814]) | ( l_39 [1569] &  i[1814]);
assign l_38[1306]    = ( l_39 [1570] & !i[1814]) | ( l_39 [1571] &  i[1814]);
assign l_38[1307]    = ( l_39 [1572] & !i[1814]) | ( l_39 [1573] &  i[1814]);
assign l_38[1308]    = ( l_39 [1574] & !i[1814]) | ( l_39 [1575] &  i[1814]);
assign l_38[1309]    = ( l_39 [1576] & !i[1814]) | ( l_39 [1577] &  i[1814]);
assign l_38[1310]    = ( l_39 [1578] & !i[1814]) | ( l_39 [1579] &  i[1814]);
assign l_38[1311]    = ( l_39 [1580] & !i[1814]) | ( l_39 [1581] &  i[1814]);
assign l_38[1312]    = ( l_39 [1582] & !i[1814]) | ( l_39 [1583] &  i[1814]);
assign l_38[1313]    = ( l_39 [1584] & !i[1814]) | ( l_39 [1585] &  i[1814]);
assign l_38[1314]    = ( l_39 [1586] & !i[1814]) | ( l_39 [1587] &  i[1814]);
assign l_38[1315]    = ( l_39 [1588] & !i[1814]) | ( l_39 [1589] &  i[1814]);
assign l_38[1316]    = ( l_39 [1590] & !i[1814]) | ( l_39 [1591] &  i[1814]);
assign l_38[1317]    = ( l_39 [1592] & !i[1814]) | ( l_39 [1593] &  i[1814]);
assign l_38[1318]    = ( l_39 [1594] & !i[1814]) | ( l_39 [1595] &  i[1814]);
assign l_38[1319]    = ( l_39 [1596] & !i[1814]) | ( l_39 [1597] &  i[1814]);
assign l_38[1320]    = ( l_39 [1598] & !i[1814]) | ( l_39 [1599] &  i[1814]);
assign l_38[1321]    = ( l_39 [1600] & !i[1814]) | ( l_39 [1601] &  i[1814]);
assign l_38[1322]    = ( l_39 [1602] & !i[1814]) | ( l_39 [1603] &  i[1814]);
assign l_38[1323]    = ( l_39 [1604] & !i[1814]) | ( l_39 [1605] &  i[1814]);
assign l_38[1324]    = ( l_39 [1606] & !i[1814]) | ( l_39 [1607] &  i[1814]);
assign l_38[1325]    = ( l_39 [1608] & !i[1814]) | ( l_39 [1609] &  i[1814]);
assign l_38[1326]    = ( l_39 [1610] & !i[1814]) | ( l_39 [1611] &  i[1814]);
assign l_38[1327]    = ( l_39 [1612] & !i[1814]) | ( l_39 [1613] &  i[1814]);
assign l_38[1328]    = ( l_39 [1614] & !i[1814]) | ( l_39 [1615] &  i[1814]);
assign l_38[1329]    = ( l_39 [1616] & !i[1814]) | ( l_39 [1617] &  i[1814]);
assign l_38[1330]    = ( l_39 [1618] & !i[1814]) | ( l_39 [1619] &  i[1814]);
assign l_38[1331]    = ( l_39 [1620] & !i[1814]) | ( l_39 [1621] &  i[1814]);
assign l_38[1332]    = ( l_39 [1622] & !i[1814]) | ( l_39 [1623] &  i[1814]);
assign l_38[1333]    = ( l_39 [1624] & !i[1814]) | ( l_39 [1625] &  i[1814]);
assign l_38[1334]    = ( l_39 [1626] & !i[1814]) | ( l_39 [1627] &  i[1814]);
assign l_38[1335]    = ( l_39 [1628] & !i[1814]) | ( l_39 [1629] &  i[1814]);
assign l_38[1336]    = ( l_39 [1630] & !i[1814]) | ( l_39 [1631] &  i[1814]);
assign l_38[1337]    = ( l_39 [1632] & !i[1814]) | ( l_39 [1633] &  i[1814]);
assign l_38[1338]    = ( l_39 [1634] & !i[1814]) | ( l_39 [1635] &  i[1814]);
assign l_38[1339]    = ( l_39 [1636] & !i[1814]) | ( l_39 [1637] &  i[1814]);
assign l_38[1340]    = ( l_39 [1638] & !i[1814]) | ( l_39 [1639] &  i[1814]);
assign l_38[1341]    = ( l_39 [1640] & !i[1814]) | ( l_39 [1641] &  i[1814]);
assign l_38[1342]    = ( l_39 [1642] & !i[1814]) | ( l_39 [1643] &  i[1814]);
assign l_38[1343]    = ( l_39 [1644] & !i[1814]) | ( l_39 [1645] &  i[1814]);
assign l_38[1344]    = ( l_39 [1646] & !i[1814]) | ( l_39 [1647] &  i[1814]);
assign l_38[1345]    = ( l_39 [1648] & !i[1814]) | ( l_39 [1649] &  i[1814]);
assign l_38[1346]    = ( l_39 [1650] & !i[1814]) | ( l_39 [1651] &  i[1814]);
assign l_38[1347]    = ( l_39 [1652] & !i[1814]) | ( l_39 [1653] &  i[1814]);
assign l_38[1348]    = ( l_39 [1654] & !i[1814]) | ( l_39 [1655] &  i[1814]);
assign l_38[1349]    = ( l_39 [1656] & !i[1814]) | ( l_39 [1657] &  i[1814]);
assign l_38[1350]    = ( l_39 [1658] & !i[1814]) | ( l_39 [1659] &  i[1814]);
assign l_38[1351]    = ( l_39 [1660] & !i[1814]) | ( l_39 [1661] &  i[1814]);
assign l_38[1352]    = ( l_39 [1662] & !i[1814]) | ( l_39 [1663] &  i[1814]);
assign l_38[1353]    = ( l_39 [1664] & !i[1814]) | ( l_39 [1665] &  i[1814]);
assign l_38[1354]    = ( l_39 [1666] & !i[1814]) | ( l_39 [1667] &  i[1814]);
assign l_38[1355]    = ( l_39 [1668] & !i[1814]) | ( l_39 [1669] &  i[1814]);
assign l_38[1356]    = ( l_39 [1670] & !i[1814]) | ( l_39 [1671] &  i[1814]);
assign l_38[1357]    = ( l_39 [1672] & !i[1814]) | ( l_39 [1673] &  i[1814]);
assign l_38[1358]    = ( l_39 [1674] & !i[1814]) | ( l_39 [1675] &  i[1814]);
assign l_38[1359]    = ( l_39 [1676] & !i[1814]) | ( l_39 [1677] &  i[1814]);
assign l_38[1360]    = ( l_39 [1678] & !i[1814]) | ( l_39 [1679] &  i[1814]);
assign l_38[1361]    = ( l_39 [1680] & !i[1814]) | ( l_39 [1681] &  i[1814]);
assign l_38[1362]    = ( l_39 [1682] & !i[1814]) | ( l_39 [1683] &  i[1814]);
assign l_38[1363]    = ( l_39 [1684] & !i[1814]) | ( l_39 [1685] &  i[1814]);
assign l_38[1364]    = ( l_39 [1686] & !i[1814]) | ( l_39 [1687] &  i[1814]);
assign l_38[1365]    = ( l_39 [1688] & !i[1814]) | ( l_39 [1689] &  i[1814]);
assign l_38[1366]    = ( l_39 [1690] & !i[1814]) | ( l_39 [1691] &  i[1814]);
assign l_38[1367]    = ( l_39 [1692] & !i[1814]) | ( l_39 [1693] &  i[1814]);
assign l_38[1368]    = ( l_39 [1694] & !i[1814]) | ( l_39 [1695] &  i[1814]);
assign l_38[1369]    = ( l_39 [1696] & !i[1814]) | ( l_39 [1697] &  i[1814]);
assign l_38[1370]    = ( l_39 [1698] & !i[1814]) | ( l_39 [1699] &  i[1814]);
assign l_38[1371]    = ( l_39 [1700] & !i[1814]) | ( l_39 [1701] &  i[1814]);
assign l_38[1372]    = ( l_39 [1702] & !i[1814]) | ( l_39 [1703] &  i[1814]);
assign l_38[1373]    = ( l_39 [1704] & !i[1814]) | ( l_39 [1705] &  i[1814]);
assign l_38[1374]    = ( l_39 [1706] & !i[1814]) | ( l_39 [1707] &  i[1814]);
assign l_38[1375]    = ( l_39 [1708] & !i[1814]) | ( l_39 [1709] &  i[1814]);
assign l_38[1376]    = ( l_39 [1710] & !i[1814]) | ( l_39 [1711] &  i[1814]);
assign l_38[1377]    = ( l_39 [1712] & !i[1814]) | ( l_39 [1713] &  i[1814]);
assign l_38[1378]    = ( l_39 [1714] & !i[1814]) | ( l_39 [1715] &  i[1814]);
assign l_38[1379]    = ( l_39 [1716] & !i[1814]) | ( l_39 [1717] &  i[1814]);
assign l_38[1380]    = ( l_39 [1718] & !i[1814]) | ( l_39 [1719] &  i[1814]);
assign l_38[1381]    = ( l_39 [1720] & !i[1814]) | ( l_39 [1721] &  i[1814]);
assign l_38[1382]    = ( l_39 [1722] & !i[1814]) | ( l_39 [1723] &  i[1814]);
assign l_38[1383]    = ( l_39 [1724] & !i[1814]) | ( l_39 [1725] &  i[1814]);
assign l_38[1384]    = ( l_39 [1726] & !i[1814]) | ( l_39 [1727] &  i[1814]);
assign l_38[1385]    = ( l_39 [1728] & !i[1814]) | ( l_39 [1729] &  i[1814]);
assign l_38[1386]    = ( l_39 [1730] & !i[1814]) | ( l_39 [1731] &  i[1814]);
assign l_38[1387]    = ( l_39 [1732] & !i[1814]) | ( l_39 [1733] &  i[1814]);
assign l_38[1388]    = ( l_39 [1734] & !i[1814]) | ( l_39 [1735] &  i[1814]);
assign l_38[1389]    = ( l_39 [1736] & !i[1814]) | ( l_39 [1737] &  i[1814]);
assign l_38[1390]    = ( l_39 [1738] & !i[1814]) | ( l_39 [1739] &  i[1814]);
assign l_38[1391]    = ( l_39 [1740] & !i[1814]) | ( l_39 [1741] &  i[1814]);
assign l_38[1392]    = ( l_39 [1742] & !i[1814]) | ( l_39 [1743] &  i[1814]);
assign l_38[1393]    = ( l_39 [1744] & !i[1814]) | ( l_39 [1745] &  i[1814]);
assign l_38[1394]    = ( l_39 [1746] & !i[1814]) | ( l_39 [1747] &  i[1814]);
assign l_38[1395]    = ( l_39 [1748] & !i[1814]) | ( l_39 [1749] &  i[1814]);
assign l_38[1396]    = ( l_39 [1750] & !i[1814]) | ( l_39 [1751] &  i[1814]);
assign l_38[1397]    = ( l_39 [1752] & !i[1814]) | ( l_39 [1753] &  i[1814]);
assign l_38[1398]    = ( l_39 [1754] & !i[1814]) | ( l_39 [1755] &  i[1814]);
assign l_38[1399]    = ( l_39 [1756] & !i[1814]) | ( l_39 [1757] &  i[1814]);
assign l_38[1400]    = ( l_39 [1758] & !i[1814]) | ( l_39 [1759] &  i[1814]);
assign l_38[1401]    = ( l_39 [1760] & !i[1814]) | ( l_39 [1761] &  i[1814]);
assign l_38[1402]    = ( l_39 [1762] & !i[1814]) | ( l_39 [1763] &  i[1814]);
assign l_38[1403]    = ( l_39 [1764] & !i[1814]) | ( l_39 [1765] &  i[1814]);
assign l_38[1404]    = ( l_39 [1766] & !i[1814]) | ( l_39 [1767] &  i[1814]);
assign l_38[1405]    = ( l_39 [1768] & !i[1814]) | ( l_39 [1769] &  i[1814]);
assign l_38[1406]    = ( l_39 [1770] & !i[1814]) | ( l_39 [1771] &  i[1814]);
assign l_38[1407]    = ( l_39 [1772] & !i[1814]) | ( l_39 [1773] &  i[1814]);
assign l_38[1408]    = ( l_39 [1774] & !i[1814]) | ( l_39 [1775] &  i[1814]);
assign l_38[1409]    = ( l_39 [1776] & !i[1814]) | ( l_39 [1777] &  i[1814]);
assign l_38[1410]    = ( l_39 [1778] & !i[1814]) | ( l_39 [1779] &  i[1814]);
assign l_38[1411]    = ( l_39 [1780] & !i[1814]) | ( l_39 [1781] &  i[1814]);
assign l_38[1412]    = ( l_39 [1782] & !i[1814]) | ( l_39 [1783] &  i[1814]);
assign l_38[1413]    = ( l_39 [1784] & !i[1814]) | ( l_39 [1785] &  i[1814]);
assign l_38[1414]    = ( l_39 [1786] & !i[1814]) | ( l_39 [1787] &  i[1814]);
assign l_38[1415]    = ( l_39 [1788] & !i[1814]) | ( l_39 [1789] &  i[1814]);
assign l_38[1416]    = ( l_39 [1790] & !i[1814]) | ( l_39 [1791] &  i[1814]);
assign l_38[1417]    = ( l_39 [1792] & !i[1814]) | ( l_39 [1793] &  i[1814]);
assign l_38[1418]    = ( l_39 [1794] & !i[1814]) | ( l_39 [1795] &  i[1814]);
assign l_38[1419]    = ( l_39 [1796] & !i[1814]) | ( l_39 [1797] &  i[1814]);
assign l_38[1420]    = ( l_39 [1798] & !i[1814]) | ( l_39 [1799] &  i[1814]);
assign l_38[1421]    = ( l_39 [1800] & !i[1814]) | ( l_39 [1801] &  i[1814]);
assign l_38[1422]    = ( l_39 [1802] & !i[1814]) | ( l_39 [1803] &  i[1814]);
assign l_38[1423]    = ( l_39 [1804] & !i[1814]) | ( l_39 [1805] &  i[1814]);
assign l_38[1424]    = ( l_39 [1806] & !i[1814]) | ( l_39 [1807] &  i[1814]);
assign l_38[1425]    = ( l_39 [1808] & !i[1814]) | ( l_39 [1809] &  i[1814]);
assign l_38[1426]    = ( l_39 [1810] & !i[1814]) | ( l_39 [1811] &  i[1814]);
assign l_38[1427]    = ( l_39 [1812] & !i[1814]) | ( l_39 [1813] &  i[1814]);
assign l_38[1428]    = ( l_39 [1814] & !i[1814]) | ( l_39 [1815] &  i[1814]);
assign l_38[1429]    = ( l_39 [1816] & !i[1814]) | ( l_39 [1817] &  i[1814]);
assign l_38[1430]    = ( l_39 [1818] & !i[1814]) | ( l_39 [1819] &  i[1814]);
assign l_38[1431]    = ( l_39 [1820] & !i[1814]) | ( l_39 [1821] &  i[1814]);
assign l_38[1432]    = ( l_39 [1822] & !i[1814]) | ( l_39 [1823] &  i[1814]);
assign l_38[1433]    = ( l_39 [1824] & !i[1814]) | ( l_39 [1825] &  i[1814]);
assign l_38[1434]    = ( l_39 [1826] & !i[1814]) | ( l_39 [1827] &  i[1814]);
assign l_38[1435]    = ( l_39 [1828] & !i[1814]) | ( l_39 [1829] &  i[1814]);
assign l_38[1436]    = ( l_39 [1830] & !i[1814]) | ( l_39 [1831] &  i[1814]);
assign l_38[1437]    = ( l_39 [1832] & !i[1814]) | ( l_39 [1833] &  i[1814]);
assign l_38[1438]    = ( l_39 [1834] & !i[1814]) | ( l_39 [1835] &  i[1814]);
assign l_38[1439]    = ( l_39 [1836] & !i[1814]) | ( l_39 [1837] &  i[1814]);
assign l_38[1440]    = ( l_39 [1838] & !i[1814]) | ( l_39 [1839] &  i[1814]);
assign l_38[1441]    = ( l_39 [1840] & !i[1814]) | ( l_39 [1841] &  i[1814]);
assign l_38[1442]    = ( l_39 [1842] & !i[1814]) | ( l_39 [1843] &  i[1814]);
assign l_38[1443]    = ( l_39 [1844] & !i[1814]) | ( l_39 [1845] &  i[1814]);
assign l_38[1444]    = ( l_39 [1846] & !i[1814]) | ( l_39 [1847] &  i[1814]);
assign l_38[1445]    = ( l_39 [1848] & !i[1814]) | ( l_39 [1849] &  i[1814]);
assign l_38[1446]    = ( l_39 [1850] & !i[1814]) | ( l_39 [1851] &  i[1814]);
assign l_38[1447]    = ( l_39 [1852] & !i[1814]) | ( l_39 [1853] &  i[1814]);
assign l_38[1448]    = ( l_39 [1854] & !i[1814]) | ( l_39 [1855] &  i[1814]);
assign l_38[1449]    = ( l_39 [1856] & !i[1814]) | ( l_39 [1857] &  i[1814]);
assign l_38[1450]    = ( l_39 [1858] & !i[1814]) | ( l_39 [1859] &  i[1814]);
assign l_38[1451]    = ( l_39 [1860] & !i[1814]) | ( l_39 [1861] &  i[1814]);
assign l_38[1452]    = ( l_39 [1862] & !i[1814]) | ( l_39 [1863] &  i[1814]);
assign l_38[1453]    = ( l_39 [1864] & !i[1814]) | ( l_39 [1865] &  i[1814]);
assign l_38[1454]    = ( l_39 [1866] & !i[1814]) | ( l_39 [1867] &  i[1814]);
assign l_38[1455]    = ( l_39 [1868] & !i[1814]) | ( l_39 [1869] &  i[1814]);
assign l_38[1456]    = ( l_39 [1870] & !i[1814]) | ( l_39 [1871] &  i[1814]);
assign l_38[1457]    = ( l_39 [1872] & !i[1814]) | ( l_39 [1873] &  i[1814]);
assign l_38[1458]    = ( l_39 [1874] & !i[1814]) | ( l_39 [1875] &  i[1814]);
assign l_38[1459]    = ( l_39 [1876] & !i[1814]) | ( l_39 [1877] &  i[1814]);
assign l_38[1460]    = ( l_39 [1878] & !i[1814]) | ( l_39 [1879] &  i[1814]);
assign l_38[1461]    = ( l_39 [1880] & !i[1814]) | ( l_39 [1881] &  i[1814]);
assign l_38[1462]    = ( l_39 [1882] & !i[1814]) | ( l_39 [1883] &  i[1814]);
assign l_38[1463]    = ( l_39 [1884] & !i[1814]) | ( l_39 [1885] &  i[1814]);
assign l_38[1464]    = ( l_39 [1886] & !i[1814]) | ( l_39 [1887] &  i[1814]);
assign l_38[1465]    = ( l_39 [1888] & !i[1814]) | ( l_39 [1889] &  i[1814]);
assign l_38[1466]    = ( l_39 [1890] & !i[1814]) | ( l_39 [1891] &  i[1814]);
assign l_38[1467]    = ( l_39 [1892] & !i[1814]) | ( l_39 [1893] &  i[1814]);
assign l_38[1468]    = ( l_39 [1894] & !i[1814]) | ( l_39 [1895] &  i[1814]);
assign l_38[1469]    = ( l_39 [1896] & !i[1814]) | ( l_39 [1897] &  i[1814]);
assign l_38[1470]    = ( l_39 [1898] & !i[1814]) | ( l_39 [1899] &  i[1814]);
assign l_38[1471]    = ( l_39 [1900] & !i[1814]) | ( l_39 [1901] &  i[1814]);
assign l_38[1472]    = ( l_39 [1902] & !i[1814]) | ( l_39 [1903] &  i[1814]);
assign l_38[1473]    = ( l_39 [1904] & !i[1814]) | ( l_39 [1905] &  i[1814]);
assign l_38[1474]    = ( l_39 [1906] & !i[1814]) | ( l_39 [1907] &  i[1814]);
assign l_38[1475]    = ( l_39 [1908] & !i[1814]) | ( l_39 [1909] &  i[1814]);
assign l_38[1476]    = ( l_39 [1910] & !i[1814]) | ( l_39 [1911] &  i[1814]);
assign l_38[1477]    = ( l_39 [1912] & !i[1814]) | ( l_39 [1913] &  i[1814]);
assign l_38[1478]    = ( l_39 [1914] & !i[1814]) | ( l_39 [1915] &  i[1814]);
assign l_38[1479]    = ( l_39 [1916] & !i[1814]) | ( l_39 [1917] &  i[1814]);
assign l_38[1480]    = ( l_39 [1918] & !i[1814]) | ( l_39 [1919] &  i[1814]);
assign l_38[1481]    = ( l_39 [1920] & !i[1814]) | ( l_39 [1921] &  i[1814]);
assign l_38[1482]    = ( l_39 [1922] & !i[1814]) | ( l_39 [1923] &  i[1814]);
assign l_38[1483]    = ( l_39 [1924] & !i[1814]) | ( l_39 [1925] &  i[1814]);
assign l_38[1484]    = ( l_39 [1926] & !i[1814]) | ( l_39 [1927] &  i[1814]);
assign l_38[1485]    = ( l_39 [1928] & !i[1814]) | ( l_39 [1929] &  i[1814]);
assign l_38[1486]    = ( l_39 [1930] & !i[1814]) | ( l_39 [1931] &  i[1814]);
assign l_38[1487]    = ( l_39 [1932] & !i[1814]) | ( l_39 [1933] &  i[1814]);
assign l_38[1488]    = ( l_39 [1934] & !i[1814]) | ( l_39 [1935] &  i[1814]);
assign l_38[1489]    = ( l_39 [1936] & !i[1814]) | ( l_39 [1937] &  i[1814]);
assign l_38[1490]    = ( l_39 [1938] & !i[1814]) | ( l_39 [1939] &  i[1814]);
assign l_38[1491]    = ( l_39 [1940] & !i[1814]) | ( l_39 [1941] &  i[1814]);
assign l_38[1492]    = ( l_39 [1942] & !i[1814]) | ( l_39 [1943] &  i[1814]);
assign l_38[1493]    = ( l_39 [1944] & !i[1814]) | ( l_39 [1945] &  i[1814]);
assign l_38[1494]    = ( l_39 [1946] & !i[1814]) | ( l_39 [1947] &  i[1814]);
assign l_38[1495]    = ( l_39 [1948] & !i[1814]) | ( l_39 [1949] &  i[1814]);
assign l_38[1496]    = ( l_39 [1950] & !i[1814]) | ( l_39 [1951] &  i[1814]);
assign l_38[1497]    = ( l_39 [1952] & !i[1814]) | ( l_39 [1953] &  i[1814]);
assign l_38[1498]    = ( l_39 [1954] & !i[1814]) | ( l_39 [1955] &  i[1814]);
assign l_38[1499]    = ( l_39 [1956] & !i[1814]) | ( l_39 [1957] &  i[1814]);
assign l_38[1500]    = ( l_39 [1958] & !i[1814]) | ( l_39 [1959] &  i[1814]);
assign l_38[1501]    = ( l_39 [1960] & !i[1814]) | ( l_39 [1961] &  i[1814]);
assign l_38[1502]    = ( l_39 [1962] & !i[1814]) | ( l_39 [1963] &  i[1814]);
assign l_38[1503]    = ( l_39 [1964] & !i[1814]) | ( l_39 [1965] &  i[1814]);
assign l_38[1504]    = ( l_39 [1966] & !i[1814]) | ( l_39 [1967] &  i[1814]);
assign l_38[1505]    = ( l_39 [1968] & !i[1814]) | ( l_39 [1969] &  i[1814]);
assign l_38[1506]    = ( l_39 [1970] & !i[1814]) | ( l_39 [1971] &  i[1814]);
assign l_38[1507]    = ( l_39 [1972] & !i[1814]) | ( l_39 [1973] &  i[1814]);
assign l_38[1508]    = ( l_39 [1974] & !i[1814]) | ( l_39 [1975] &  i[1814]);
assign l_38[1509]    = ( l_39 [1976] & !i[1814]) | ( l_39 [1977] &  i[1814]);
assign l_38[1510]    = ( l_39 [1978] & !i[1814]) | ( l_39 [1979] &  i[1814]);
assign l_38[1511]    = ( l_39 [1980] & !i[1814]) | ( l_39 [1981] &  i[1814]);
assign l_38[1512]    = ( l_39 [1982] & !i[1814]) | ( l_39 [1983] &  i[1814]);
assign l_38[1513]    = ( l_39 [1984] & !i[1814]) | ( l_39 [1985] &  i[1814]);
assign l_38[1514]    = ( l_39 [1986] & !i[1814]) | ( l_39 [1987] &  i[1814]);
assign l_38[1515]    = ( l_39 [1988] & !i[1814]) | ( l_39 [1989] &  i[1814]);
assign l_38[1516]    = ( l_39 [1990] & !i[1814]) | ( l_39 [1991] &  i[1814]);
assign l_38[1517]    = ( l_39 [1992] & !i[1814]) | ( l_39 [1993] &  i[1814]);
assign l_38[1518]    = ( l_39 [1994] & !i[1814]) | ( l_39 [1995] &  i[1814]);
assign l_38[1519]    = ( l_39 [1996] & !i[1814]) | ( l_39 [1997] &  i[1814]);
assign l_38[1520]    = ( l_39 [1998] & !i[1814]) | ( l_39 [1999] &  i[1814]);
assign l_38[1521]    = ( l_39 [2000] & !i[1814]) | ( l_39 [2001] &  i[1814]);
assign l_38[1522]    = ( l_39 [2002] & !i[1814]) | ( l_39 [2003] &  i[1814]);
assign l_38[1523]    = ( l_39 [2004] & !i[1814]) | ( l_39 [2005] &  i[1814]);
assign l_38[1524]    = ( l_39 [2006] & !i[1814]) | ( l_39 [2007] &  i[1814]);
assign l_38[1525]    = ( l_39 [2008] & !i[1814]) | ( l_39 [2009] &  i[1814]);
assign l_38[1526]    = ( l_39 [2010] & !i[1814]) | ( l_39 [2011] &  i[1814]);
assign l_38[1527]    = ( l_39 [2012] & !i[1814]) | ( l_39 [2013] &  i[1814]);
assign l_38[1528]    = ( l_39 [2014] & !i[1814]) | ( l_39 [2015] &  i[1814]);
assign l_38[1529]    = ( l_39 [2016] & !i[1814]) | ( l_39 [2017] &  i[1814]);
assign l_38[1530]    = ( l_39 [2018] & !i[1814]) | ( l_39 [2019] &  i[1814]);
assign l_38[1531]    = ( l_39 [2020] & !i[1814]) | ( l_39 [2021] &  i[1814]);
assign l_38[1532]    = ( l_39 [2022] & !i[1814]) | ( l_39 [2023] &  i[1814]);
assign l_38[1533]    = ( l_39 [2024] & !i[1814]) | ( l_39 [2025] &  i[1814]);
assign l_38[1534]    = ( l_39 [2026] & !i[1814]) | ( l_39 [2027] &  i[1814]);
assign l_38[1535]    = ( l_39 [2028] & !i[1814]) | ( l_39 [2029] &  i[1814]);
assign l_38[1536]    = ( l_39 [2030] & !i[1814]) | ( l_39 [2031] &  i[1814]);
assign l_38[1537]    = ( l_39 [2032] & !i[1814]) | ( l_39 [2033] &  i[1814]);
assign l_38[1538]    = ( l_39 [2034] & !i[1814]) | ( l_39 [2035] &  i[1814]);
assign l_38[1539]    = ( l_39 [2036] & !i[1814]) | ( l_39 [2037] &  i[1814]);
assign l_38[1540]    = ( l_39 [2038] & !i[1814]) | ( l_39 [2039] &  i[1814]);
assign l_38[1541]    = ( l_39 [2040] & !i[1814]) | ( l_39 [2041] &  i[1814]);
assign l_38[1542]    = ( l_39 [2042] & !i[1814]) | ( l_39 [2043] &  i[1814]);
assign l_38[1543]    = ( l_39 [2044] & !i[1814]) | ( l_39 [2045] &  i[1814]);
assign l_38[1544]    = ( l_39 [2046] & !i[1814]) | ( l_39 [2047] &  i[1814]);
assign l_38[1545]    = ( l_39 [2048] & !i[1814]) | ( l_39 [2049] &  i[1814]);
assign l_38[1546]    = ( l_39 [2050] & !i[1814]) | ( l_39 [2051] &  i[1814]);
assign l_38[1547]    = ( l_39 [2052] & !i[1814]) | ( l_39 [2053] &  i[1814]);
assign l_38[1548]    = ( l_39 [2054] & !i[1814]) | ( l_39 [2055] &  i[1814]);
assign l_38[1549]    = ( l_39 [2056] & !i[1814]) | ( l_39 [2057] &  i[1814]);
assign l_38[1550]    = ( l_39 [2058] & !i[1814]) | ( l_39 [2059] &  i[1814]);
assign l_38[1551]    = ( l_39 [2060] & !i[1814]) | ( l_39 [2061] &  i[1814]);
assign l_38[1552]    = ( l_39 [2062] & !i[1814]) | ( l_39 [2063] &  i[1814]);
assign l_38[1553]    = ( l_39 [2064] & !i[1814]) | ( l_39 [2065] &  i[1814]);
assign l_38[1554]    = ( l_39 [2066] & !i[1814]) | ( l_39 [2067] &  i[1814]);
assign l_38[1555]    = ( l_39 [2068] & !i[1814]) | ( l_39 [2069] &  i[1814]);
assign l_38[1556]    = ( l_39 [2070] & !i[1814]) | ( l_39 [2071] &  i[1814]);
assign l_38[1557]    = ( l_39 [2072] & !i[1814]) | ( l_39 [2073] &  i[1814]);
assign l_38[1558]    = ( l_39 [2074] & !i[1814]) | ( l_39 [2075] &  i[1814]);
assign l_38[1559]    = ( l_39 [2076] & !i[1814]) | ( l_39 [2077] &  i[1814]);
assign l_38[1560]    = ( l_39 [2078] & !i[1814]) | ( l_39 [2079] &  i[1814]);
assign l_38[1561]    = ( l_39 [2080] & !i[1814]) | ( l_39 [2081] &  i[1814]);
assign l_38[1562]    = ( l_39 [2082] & !i[1814]) | ( l_39 [2083] &  i[1814]);
assign l_38[1563]    = ( l_39 [2084] & !i[1814]) | ( l_39 [2085] &  i[1814]);
assign l_38[1564]    = ( l_39 [2086] & !i[1814]) | ( l_39 [2087] &  i[1814]);
assign l_38[1565]    = ( l_39 [2088] & !i[1814]) | ( l_39 [2089] &  i[1814]);
assign l_38[1566]    = ( l_39 [2090] & !i[1814]) | ( l_39 [2091] &  i[1814]);
assign l_38[1567]    = ( l_39 [2092] & !i[1814]) | ( l_39 [2093] &  i[1814]);
assign l_38[1568]    = ( l_39 [2094] & !i[1814]) | ( l_39 [2095] &  i[1814]);
assign l_38[1569]    = ( l_39 [2096] & !i[1814]) | ( l_39 [2097] &  i[1814]);
assign l_38[1570]    = ( l_39 [2098] & !i[1814]) | ( l_39 [2099] &  i[1814]);
assign l_38[1571]    = ( l_39 [2100] & !i[1814]) | ( l_39 [2101] &  i[1814]);
assign l_38[1572]    = ( l_39 [2102] & !i[1814]) | ( l_39 [2103] &  i[1814]);
assign l_38[1573]    = ( l_39 [2104] & !i[1814]) | ( l_39 [2105] &  i[1814]);
assign l_38[1574]    = ( l_39 [2106] & !i[1814]) | ( l_39 [2107] &  i[1814]);
assign l_38[1575]    = ( l_39 [2108] & !i[1814]) | ( l_39 [2109] &  i[1814]);
assign l_38[1576]    = ( l_39 [2110] & !i[1814]) | ( l_39 [2111] &  i[1814]);
assign l_38[1577]    = ( l_39 [2112] & !i[1814]) | ( l_39 [2113] &  i[1814]);
assign l_38[1578]    = ( l_39 [2114] & !i[1814]) | ( l_39 [2115] &  i[1814]);
assign l_38[1579]    = ( l_39 [2116] & !i[1814]) | ( l_39 [2117] &  i[1814]);
assign l_38[1580]    = ( l_39 [2118] & !i[1814]) | ( l_39 [2119] &  i[1814]);
assign l_38[1581]    = ( l_39 [2120] & !i[1814]) | ( l_39 [2121] &  i[1814]);
assign l_38[1582]    = ( l_39 [2122] & !i[1814]) | ( l_39 [2123] &  i[1814]);
assign l_38[1583]    = ( l_39 [2124] & !i[1814]) | ( l_39 [2125] &  i[1814]);
assign l_38[1584]    = ( l_39 [2126] & !i[1814]) | ( l_39 [2127] &  i[1814]);
assign l_38[1585]    = ( l_39 [2128] & !i[1814]) | ( l_39 [2129] &  i[1814]);
assign l_38[1586]    = ( l_39 [2130] & !i[1814]) | ( l_39 [2131] &  i[1814]);
assign l_38[1587]    = ( l_39 [2132] & !i[1814]) | ( l_39 [2133] &  i[1814]);
assign l_38[1588]    = ( l_39 [2134] & !i[1814]) | ( l_39 [2135] &  i[1814]);
assign l_38[1589]    = ( l_39 [2136] & !i[1814]) | ( l_39 [2137] &  i[1814]);
assign l_38[1590]    = ( l_39 [2138] & !i[1814]) | ( l_39 [2139] &  i[1814]);
assign l_38[1591]    = ( l_39 [2140] & !i[1814]) | ( l_39 [2141] &  i[1814]);
assign l_38[1592]    = ( l_39 [2142] & !i[1814]) | ( l_39 [2143] &  i[1814]);
assign l_38[1593]    = ( l_39 [2144] & !i[1814]) | ( l_39 [2145] &  i[1814]);
assign l_38[1594]    = ( l_39 [2146] & !i[1814]) | ( l_39 [2147] &  i[1814]);
assign l_38[1595]    = ( l_39 [2148] & !i[1814]) | ( l_39 [2149] &  i[1814]);
assign l_38[1596]    = ( l_39 [2150] & !i[1814]) | ( l_39 [2151] &  i[1814]);
assign l_38[1597]    = ( l_39 [2152] & !i[1814]) | ( l_39 [2153] &  i[1814]);
assign l_38[1598]    = ( l_39 [2154] & !i[1814]) | ( l_39 [2155] &  i[1814]);
assign l_38[1599]    = ( l_39 [2156] & !i[1814]) | ( l_39 [2157] &  i[1814]);
assign l_38[1600]    = ( l_39 [2158] & !i[1814]) | ( l_39 [2159] &  i[1814]);
assign l_38[1601]    = ( l_39 [2160] & !i[1814]) | ( l_39 [2161] &  i[1814]);
assign l_38[1602]    = ( l_39 [2162] & !i[1814]) | ( l_39 [2163] &  i[1814]);
assign l_38[1603]    = ( l_39 [2164] & !i[1814]) | ( l_39 [2165] &  i[1814]);
assign l_38[1604]    = ( l_39 [2166] & !i[1814]) | ( l_39 [2167] &  i[1814]);
assign l_38[1605]    = ( l_39 [2168] & !i[1814]) | ( l_39 [2169] &  i[1814]);
assign l_38[1606]    = ( l_39 [2170] & !i[1814]) | ( l_39 [2171] &  i[1814]);
assign l_38[1607]    = ( l_39 [2172] & !i[1814]) | ( l_39 [2173] &  i[1814]);
assign l_38[1608]    = ( l_39 [2174] & !i[1814]) | ( l_39 [2175] &  i[1814]);
assign l_38[1609]    = ( l_39 [2176] & !i[1814]) | ( l_39 [2177] &  i[1814]);
assign l_38[1610]    = ( l_39 [2178] & !i[1814]) | ( l_39 [2179] &  i[1814]);
assign l_38[1611]    = ( l_39 [2180] & !i[1814]) | ( l_39 [2181] &  i[1814]);
assign l_38[1612]    = ( l_39 [2182] & !i[1814]) | ( l_39 [2183] &  i[1814]);
assign l_38[1613]    = ( l_39 [2184] & !i[1814]) | ( l_39 [2185] &  i[1814]);
assign l_38[1614]    = ( l_39 [2186] & !i[1814]) | ( l_39 [2187] &  i[1814]);
assign l_38[1615]    = ( l_39 [2188] & !i[1814]) | ( l_39 [2189] &  i[1814]);
assign l_38[1616]    = ( l_39 [2190] & !i[1814]) | ( l_39 [2191] &  i[1814]);
assign l_38[1617]    = ( l_39 [2192] & !i[1814]) | ( l_39 [2193] &  i[1814]);
assign l_38[1618]    = ( l_39 [2194] & !i[1814]) | ( l_39 [2195] &  i[1814]);
assign l_38[1619]    = ( l_39 [2196] & !i[1814]) | ( l_39 [2197] &  i[1814]);
assign l_38[1620]    = ( l_39 [2198] & !i[1814]) | ( l_39 [2199] &  i[1814]);
assign l_38[1621]    = ( l_39 [2200] & !i[1814]) | ( l_39 [2201] &  i[1814]);
assign l_38[1622]    = ( l_39 [2202] & !i[1814]) | ( l_39 [2203] &  i[1814]);
assign l_38[1623]    = ( l_39 [2204] & !i[1814]) | ( l_39 [2205] &  i[1814]);
assign l_38[1624]    = ( l_39 [2206] & !i[1814]) | ( l_39 [2207] &  i[1814]);
assign l_38[1625]    = ( l_39 [2208] & !i[1814]) | ( l_39 [2209] &  i[1814]);
assign l_38[1626]    = ( l_39 [2210] & !i[1814]) | ( l_39 [2211] &  i[1814]);
assign l_38[1627]    = ( l_39 [2212] & !i[1814]) | ( l_39 [2213] &  i[1814]);
assign l_38[1628]    = ( l_39 [2214] & !i[1814]) | ( l_39 [2215] &  i[1814]);
assign l_38[1629]    = ( l_39 [2216] & !i[1814]) | ( l_39 [2217] &  i[1814]);
assign l_38[1630]    = ( l_39 [2218] & !i[1814]) | ( l_39 [2219] &  i[1814]);
assign l_38[1631]    = ( l_39 [2220] & !i[1814]) | ( l_39 [2221] &  i[1814]);
assign l_38[1632]    = ( l_39 [2222] & !i[1814]) | ( l_39 [2223] &  i[1814]);
assign l_38[1633]    = ( l_39 [2224] & !i[1814]) | ( l_39 [2225] &  i[1814]);
assign l_38[1634]    = ( l_39 [2226] & !i[1814]) | ( l_39 [2227] &  i[1814]);
assign l_38[1635]    = ( l_39 [2228] & !i[1814]) | ( l_39 [2229] &  i[1814]);
assign l_38[1636]    = ( l_39 [2230] & !i[1814]) | ( l_39 [2231] &  i[1814]);
assign l_38[1637]    = ( l_39 [2232] & !i[1814]) | ( l_39 [2233] &  i[1814]);
assign l_38[1638]    = ( l_39 [2234] & !i[1814]) | ( l_39 [2235] &  i[1814]);
assign l_38[1639]    = ( l_39 [2236] & !i[1814]) | ( l_39 [2237] &  i[1814]);
assign l_38[1640]    = ( l_39 [2238] & !i[1814]) | ( l_39 [2239] &  i[1814]);
assign l_38[1641]    = ( l_39 [2240] & !i[1814]) | ( l_39 [2241] &  i[1814]);
assign l_38[1642]    = ( l_39 [2242] & !i[1814]) | ( l_39 [2243] &  i[1814]);
assign l_38[1643]    = ( l_39 [2244] & !i[1814]) | ( l_39 [2245] &  i[1814]);
assign l_38[1644]    = ( l_39 [2246] & !i[1814]) | ( l_39 [2247] &  i[1814]);
assign l_38[1645]    = ( l_39 [2248] & !i[1814]) | ( l_39 [2249] &  i[1814]);
assign l_38[1646]    = ( l_39 [2250] & !i[1814]) | ( l_39 [2251] &  i[1814]);
assign l_38[1647]    = ( l_39 [2252] & !i[1814]) | ( l_39 [2253] &  i[1814]);
assign l_38[1648]    = ( l_39 [2254] & !i[1814]) | ( l_39 [2255] &  i[1814]);
assign l_38[1649]    = ( l_39 [2256] & !i[1814]) | ( l_39 [2257] &  i[1814]);
assign l_38[1650]    = ( l_39 [2258] & !i[1814]) | ( l_39 [2259] &  i[1814]);
assign l_38[1651]    = ( l_39 [2260] & !i[1814]) | ( l_39 [2261] &  i[1814]);
assign l_38[1652]    = ( l_39 [2262] & !i[1814]) | ( l_39 [2263] &  i[1814]);
assign l_38[1653]    = ( l_39 [2264] & !i[1814]) | ( l_39 [2265] &  i[1814]);
assign l_38[1654]    = ( l_39 [2266] & !i[1814]) | ( l_39 [2267] &  i[1814]);
assign l_38[1655]    = ( l_39 [2268] & !i[1814]) | ( l_39 [2269] &  i[1814]);
assign l_38[1656]    = ( l_39 [2270] & !i[1814]) | ( l_39 [2271] &  i[1814]);
assign l_38[1657]    = ( l_39 [2272] & !i[1814]) | ( l_39 [2273] &  i[1814]);
assign l_38[1658]    = ( l_39 [2274] & !i[1814]) | ( l_39 [2275] &  i[1814]);
assign l_38[1659]    = ( l_39 [2276] & !i[1814]) | ( l_39 [2277] &  i[1814]);
assign l_38[1660]    = ( l_39 [2278] & !i[1814]) | ( l_39 [2279] &  i[1814]);
assign l_38[1661]    = ( l_39 [2280] & !i[1814]) | ( l_39 [2281] &  i[1814]);
assign l_38[1662]    = ( l_39 [2282] & !i[1814]) | ( l_39 [2283] &  i[1814]);
assign l_38[1663]    = ( l_39 [2284] & !i[1814]) | ( l_39 [2285] &  i[1814]);
assign l_38[1664]    = ( l_39 [2286] & !i[1814]) | ( l_39 [2287] &  i[1814]);
assign l_38[1665]    = ( l_39 [2288] & !i[1814]) | ( l_39 [2289] &  i[1814]);
assign l_38[1666]    = ( l_39 [2290] & !i[1814]) | ( l_39 [2291] &  i[1814]);
assign l_38[1667]    = ( l_39 [2292] & !i[1814]) | ( l_39 [2293] &  i[1814]);
assign l_38[1668]    = ( l_39 [2294] & !i[1814]) | ( l_39 [2295] &  i[1814]);
assign l_38[1669]    = ( l_39 [2296] & !i[1814]) | ( l_39 [2297] &  i[1814]);
assign l_38[1670]    = ( l_39 [2298] & !i[1814]) | ( l_39 [2299] &  i[1814]);
assign l_38[1671]    = ( l_39 [2300] & !i[1814]) | ( l_39 [2301] &  i[1814]);
assign l_38[1672]    = ( l_39 [2302] & !i[1814]) | ( l_39 [2303] &  i[1814]);
assign l_38[1673]    = ( l_39 [2304] & !i[1814]) | ( l_39 [2305] &  i[1814]);
assign l_38[1674]    = ( l_39 [2306] & !i[1814]) | ( l_39 [2307] &  i[1814]);
assign l_38[1675]    = ( l_39 [2308] & !i[1814]) | ( l_39 [2309] &  i[1814]);
assign l_38[1676]    = ( l_39 [2310] & !i[1814]) | ( l_39 [2311] &  i[1814]);
assign l_38[1677]    = ( l_39 [2312] & !i[1814]) | ( l_39 [2313] &  i[1814]);
assign l_38[1678]    = ( l_39 [2314] & !i[1814]) | ( l_39 [2315] &  i[1814]);
assign l_38[1679]    = ( l_39 [2316] & !i[1814]) | ( l_39 [2317] &  i[1814]);
assign l_38[1680]    = ( l_39 [2318] & !i[1814]) | ( l_39 [2319] &  i[1814]);
assign l_38[1681]    = ( l_39 [2320] & !i[1814]) | ( l_39 [2321] &  i[1814]);
assign l_38[1682]    = ( l_39 [2322] & !i[1814]) | ( l_39 [2323] &  i[1814]);
assign l_38[1683]    = ( l_39 [2324] & !i[1814]) | ( l_39 [2325] &  i[1814]);
assign l_38[1684]    = ( l_39 [2326] & !i[1814]) | ( l_39 [2327] &  i[1814]);
assign l_38[1685]    = ( l_39 [2328] & !i[1814]) | ( l_39 [2329] &  i[1814]);
assign l_38[1686]    = ( l_39 [2330] & !i[1814]) | ( l_39 [2331] &  i[1814]);
assign l_38[1687]    = ( l_39 [2332] & !i[1814]) | ( l_39 [2333] &  i[1814]);
assign l_38[1688]    = ( l_39 [2334] & !i[1814]) | ( l_39 [2335] &  i[1814]);
assign l_38[1689]    = ( l_39 [2336] & !i[1814]) | ( l_39 [2337] &  i[1814]);
assign l_38[1690]    = ( l_39 [2338] & !i[1814]) | ( l_39 [2339] &  i[1814]);
assign l_38[1691]    = ( l_39 [2340] & !i[1814]) | ( l_39 [2341] &  i[1814]);
assign l_38[1692]    = ( l_39 [2342] & !i[1814]) | ( l_39 [2343] &  i[1814]);
assign l_38[1693]    = ( l_39 [2344] & !i[1814]) | ( l_39 [2345] &  i[1814]);
assign l_38[1694]    = ( l_39 [2346] & !i[1814]) | ( l_39 [2347] &  i[1814]);
assign l_38[1695]    = ( l_39 [2348] & !i[1814]) | ( l_39 [2349] &  i[1814]);
assign l_38[1696]    = ( l_39 [2350] & !i[1814]) | ( l_39 [2351] &  i[1814]);
assign l_38[1697]    = ( l_39 [2352] & !i[1814]) | ( l_39 [2353] &  i[1814]);
assign l_38[1698]    = ( l_39 [2354] & !i[1814]) | ( l_39 [2355] &  i[1814]);
assign l_38[1699]    = ( l_39 [2356] & !i[1814]) | ( l_39 [2357] &  i[1814]);
assign l_38[1700]    = ( l_39 [2358] & !i[1814]) | ( l_39 [2359] &  i[1814]);
assign l_38[1701]    = ( l_39 [2360] & !i[1814]) | ( l_39 [2361] &  i[1814]);
assign l_38[1702]    = ( l_39 [2362] & !i[1814]) | ( l_39 [2363] &  i[1814]);
assign l_38[1703]    = ( l_39 [2364] & !i[1814]) | ( l_39 [2365] &  i[1814]);
assign l_38[1704]    = ( l_39 [2366] & !i[1814]) | ( l_39 [2367] &  i[1814]);
assign l_38[1705]    = ( l_39 [2368] & !i[1814]) | ( l_39 [2369] &  i[1814]);
assign l_38[1706]    = ( l_39 [2370] & !i[1814]) | ( l_39 [2371] &  i[1814]);
assign l_38[1707]    = ( l_39 [2372] & !i[1814]) | ( l_39 [2373] &  i[1814]);
assign l_38[1708]    = ( l_39 [2374] & !i[1814]) | ( l_39 [2375] &  i[1814]);
assign l_38[1709]    = ( l_39 [2376] & !i[1814]) | ( l_39 [2377] &  i[1814]);
assign l_38[1710]    = ( l_39 [2378] & !i[1814]) | ( l_39 [2379] &  i[1814]);
assign l_38[1711]    = ( l_39 [2380] & !i[1814]) | ( l_39 [2381] &  i[1814]);
assign l_38[1712]    = ( l_39 [2382] & !i[1814]) | ( l_39 [2383] &  i[1814]);
assign l_38[1713]    = ( l_39 [2384] & !i[1814]) | ( l_39 [2385] &  i[1814]);
assign l_38[1714]    = ( l_39 [2386] & !i[1814]) | ( l_39 [2387] &  i[1814]);
assign l_38[1715]    = ( l_39 [2388] & !i[1814]) | ( l_39 [2389] &  i[1814]);
assign l_38[1716]    = ( l_39 [2390] & !i[1814]) | ( l_39 [2391] &  i[1814]);
assign l_38[1717]    = ( l_39 [2392] & !i[1814]) | ( l_39 [2393] &  i[1814]);
assign l_38[1718]    = ( l_39 [2394] & !i[1814]) | ( l_39 [2395] &  i[1814]);
assign l_38[1719]    = ( l_39 [2396] & !i[1814]) | ( l_39 [2397] &  i[1814]);
assign l_38[1720]    = ( l_39 [2398] & !i[1814]) | ( l_39 [2399] &  i[1814]);
assign l_38[1721]    = ( l_39 [2400] & !i[1814]) | ( l_39 [2401] &  i[1814]);
assign l_38[1722]    = ( l_39 [2402] & !i[1814]) | ( l_39 [2403] &  i[1814]);
assign l_38[1723]    = ( l_39 [2404] & !i[1814]) | ( l_39 [2405] &  i[1814]);
assign l_38[1724]    = ( l_39 [2406] & !i[1814]) | ( l_39 [2407] &  i[1814]);
assign l_38[1725]    = ( l_39 [2408] & !i[1814]) | ( l_39 [2409] &  i[1814]);
assign l_38[1726]    = ( l_39 [2410] & !i[1814]) | ( l_39 [2411] &  i[1814]);
assign l_38[1727]    = ( l_39 [2412] & !i[1814]) | ( l_39 [2413] &  i[1814]);
assign l_38[1728]    = ( l_39 [2414] & !i[1814]) | ( l_39 [2415] &  i[1814]);
assign l_38[1729]    = ( l_39 [2416] & !i[1814]) | ( l_39 [2417] &  i[1814]);
assign l_38[1730]    = ( l_39 [2418] & !i[1814]) | ( l_39 [2419] &  i[1814]);
assign l_38[1731]    = ( l_39 [2420] & !i[1814]) | ( l_39 [2421] &  i[1814]);
assign l_38[1732]    = ( l_39 [2422] & !i[1814]) | ( l_39 [2423] &  i[1814]);
assign l_38[1733]    = ( l_39 [2424] & !i[1814]) | ( l_39 [2425] &  i[1814]);
assign l_38[1734]    = ( l_39 [2426] & !i[1814]) | ( l_39 [2427] &  i[1814]);
assign l_38[1735]    = ( l_39 [2428] & !i[1814]) | ( l_39 [2429] &  i[1814]);
assign l_38[1736]    = ( l_39 [2430] & !i[1814]) | ( l_39 [2431] &  i[1814]);
assign l_38[1737]    = ( l_39 [2432] & !i[1814]) | ( l_39 [2433] &  i[1814]);
assign l_38[1738]    = ( l_39 [2434] & !i[1814]) | ( l_39 [2435] &  i[1814]);
assign l_38[1739]    = ( l_39 [2436] & !i[1814]) | ( l_39 [2437] &  i[1814]);
assign l_38[1740]    = ( l_39 [2438] & !i[1814]) | ( l_39 [2439] &  i[1814]);
assign l_38[1741]    = ( l_39 [2440] & !i[1814]) | ( l_39 [2441] &  i[1814]);
assign l_38[1742]    = ( l_39 [2442] & !i[1814]) | ( l_39 [2443] &  i[1814]);
assign l_38[1743]    = ( l_39 [2444] & !i[1814]) | ( l_39 [2445] &  i[1814]);
assign l_38[1744]    = ( l_39 [2446] & !i[1814]) | ( l_39 [2447] &  i[1814]);
assign l_38[1745]    = ( l_39 [2448] & !i[1814]) | ( l_39 [2449] &  i[1814]);
assign l_38[1746]    = ( l_39 [2450] & !i[1814]) | ( l_39 [2451] &  i[1814]);
assign l_38[1747]    = ( l_39 [2452] & !i[1814]) | ( l_39 [2453] &  i[1814]);
assign l_38[1748]    = ( l_39 [2454] & !i[1814]) | ( l_39 [2455] &  i[1814]);
assign l_38[1749]    = ( l_39 [2456] & !i[1814]) | ( l_39 [2457] &  i[1814]);
assign l_38[1750]    = ( l_39 [2458] & !i[1814]) | ( l_39 [2459] &  i[1814]);
assign l_38[1751]    = ( l_39 [2460] & !i[1814]) | ( l_39 [2461] &  i[1814]);
assign l_38[1752]    = ( l_39 [2462] & !i[1814]) | ( l_39 [2463] &  i[1814]);
assign l_38[1753]    = ( l_39 [2464] & !i[1814]) | ( l_39 [2465] &  i[1814]);
assign l_38[1754]    = ( l_39 [2466] & !i[1814]) | ( l_39 [2467] &  i[1814]);
assign l_38[1755]    = ( l_39 [2468] & !i[1814]) | ( l_39 [2469] &  i[1814]);
assign l_38[1756]    = ( l_39 [2470] & !i[1814]) | ( l_39 [2471] &  i[1814]);
assign l_38[1757]    = ( l_39 [2472] & !i[1814]) | ( l_39 [2473] &  i[1814]);
assign l_38[1758]    = ( l_39 [2474] & !i[1814]) | ( l_39 [2475] &  i[1814]);
assign l_38[1759]    = ( l_39 [2476] & !i[1814]) | ( l_39 [2477] &  i[1814]);
assign l_38[1760]    = ( l_39 [2478] & !i[1814]) | ( l_39 [2479] &  i[1814]);
assign l_38[1761]    = ( l_39 [2480] & !i[1814]) | ( l_39 [2481] &  i[1814]);
assign l_38[1762]    = ( l_39 [2482] & !i[1814]) | ( l_39 [2483] &  i[1814]);
assign l_38[1763]    = ( l_39 [2484] & !i[1814]) | ( l_39 [2485] &  i[1814]);
assign l_38[1764]    = ( l_39 [2486] & !i[1814]) | ( l_39 [2487] &  i[1814]);
assign l_38[1765]    = ( l_39 [2488] & !i[1814]) | ( l_39 [2489] &  i[1814]);
assign l_38[1766]    = ( l_39 [2490] & !i[1814]) | ( l_39 [2491] &  i[1814]);
assign l_38[1767]    = ( l_39 [2492] & !i[1814]) | ( l_39 [2493] &  i[1814]);
assign l_38[1768]    = ( l_39 [2494] & !i[1814]) | ( l_39 [2495] &  i[1814]);
assign l_38[1769]    = ( l_39 [2496] & !i[1814]) | ( l_39 [2497] &  i[1814]);
assign l_38[1770]    = ( l_39 [2498] & !i[1814]) | ( l_39 [2499] &  i[1814]);
assign l_38[1771]    = ( l_39 [2500] & !i[1814]) | ( l_39 [2501] &  i[1814]);
assign l_38[1772]    = ( l_39 [2502] & !i[1814]) | ( l_39 [2503] &  i[1814]);
assign l_38[1773]    = ( l_39 [2504] & !i[1814]) | ( l_39 [2505] &  i[1814]);
assign l_38[1774]    = ( l_39 [2506] & !i[1814]) | ( l_39 [2507] &  i[1814]);
assign l_38[1775]    = ( l_39 [2508] & !i[1814]) | ( l_39 [2509] &  i[1814]);
assign l_38[1776]    = ( l_39 [2510] & !i[1814]) | ( l_39 [2511] &  i[1814]);
assign l_38[1777]    = ( l_39 [2512] & !i[1814]) | ( l_39 [2513] &  i[1814]);
assign l_38[1778]    = ( l_39 [2514] & !i[1814]) | ( l_39 [2515] &  i[1814]);
assign l_38[1779]    = ( l_39 [2516] & !i[1814]) | ( l_39 [2517] &  i[1814]);
assign l_38[1780]    = ( l_39 [2518] & !i[1814]) | ( l_39 [2519] &  i[1814]);
assign l_38[1781]    = ( l_39 [2520] & !i[1814]) | ( l_39 [2521] &  i[1814]);
assign l_38[1782]    = ( l_39 [2522] & !i[1814]) | ( l_39 [2523] &  i[1814]);
assign l_38[1783]    = ( l_39 [2524] & !i[1814]) | ( l_39 [2525] &  i[1814]);
assign l_38[1784]    = ( l_39 [2526] & !i[1814]) | ( l_39 [2527] &  i[1814]);
assign l_38[1785]    = ( l_39 [2528] & !i[1814]) | ( l_39 [2529] &  i[1814]);
assign l_38[1786]    = ( l_39 [2530] & !i[1814]) | ( l_39 [2531] &  i[1814]);
assign l_38[1787]    = ( l_39 [2532] & !i[1814]) | ( l_39 [2533] &  i[1814]);
assign l_38[1788]    = ( l_39 [2534] & !i[1814]) | ( l_39 [2535] &  i[1814]);
assign l_38[1789]    = ( l_39 [2536] & !i[1814]) | ( l_39 [2537] &  i[1814]);
assign l_38[1790]    = ( l_39 [2538] & !i[1814]) | ( l_39 [2539] &  i[1814]);
assign l_38[1791]    = ( l_39 [2540] & !i[1814]) | ( l_39 [2541] &  i[1814]);
assign l_38[1792]    = ( l_39 [2542] & !i[1814]) | ( l_39 [2543] &  i[1814]);
assign l_38[1793]    = ( l_39 [2544] & !i[1814]) | ( l_39 [2545] &  i[1814]);
assign l_38[1794]    = ( l_39 [2546] & !i[1814]) | ( l_39 [2547] &  i[1814]);
assign l_38[1795]    = ( l_39 [2548] & !i[1814]) | ( l_39 [2549] &  i[1814]);
assign l_38[1796]    = ( l_39 [2550] & !i[1814]) | ( l_39 [2551] &  i[1814]);
assign l_38[1797]    = ( l_39 [2552] & !i[1814]) | ( l_39 [2553] &  i[1814]);
assign l_38[1798]    = ( l_39 [2554] & !i[1814]) | ( l_39 [2555] &  i[1814]);
assign l_38[1799]    = ( l_39 [2556] & !i[1814]) | ( l_39 [2557] &  i[1814]);
assign l_38[1800]    = ( l_39 [2558] & !i[1814]) | ( l_39 [2559] &  i[1814]);
assign l_38[1801]    = ( l_39 [2560] & !i[1814]) | ( l_39 [2561] &  i[1814]);
assign l_38[1802]    = ( l_39 [2562] & !i[1814]) | ( l_39 [2563] &  i[1814]);
assign l_38[1803]    = ( l_39 [2564] & !i[1814]) | ( l_39 [2565] &  i[1814]);
assign l_38[1804]    = ( l_39 [2566] & !i[1814]) | ( l_39 [2567] &  i[1814]);
assign l_38[1805]    = ( l_39 [2568] & !i[1814]) | ( l_39 [2569] &  i[1814]);
assign l_38[1806]    = ( l_39 [2570] & !i[1814]) | ( l_39 [2571] &  i[1814]);
assign l_38[1807]    = ( l_39 [2572] & !i[1814]) | ( l_39 [2573] &  i[1814]);
assign l_38[1808]    = ( l_39 [2574] & !i[1814]) | ( l_39 [2575] &  i[1814]);
assign l_38[1809]    = ( l_39 [2576] & !i[1814]) | ( l_39 [2577] &  i[1814]);
assign l_38[1810]    = ( l_39 [2578] & !i[1814]) | ( l_39 [2579] &  i[1814]);
assign l_38[1811]    = ( l_39 [2580] & !i[1814]) | ( l_39 [2581] &  i[1814]);
assign l_38[1812]    = ( l_39 [2582] & !i[1814]) | ( l_39 [2583] &  i[1814]);
assign l_38[1813]    = ( l_39 [2584] & !i[1814]) | ( l_39 [2585] &  i[1814]);
assign l_38[1814]    = ( l_39 [2586] & !i[1814]) | ( l_39 [2587] &  i[1814]);
assign l_38[1815]    = ( l_39 [2588] & !i[1814]) | ( l_39 [2589] &  i[1814]);
assign l_38[1816]    = ( l_39 [2590] & !i[1814]) | ( l_39 [2591] &  i[1814]);
assign l_38[1817]    = ( l_39 [2592] & !i[1814]) | ( l_39 [2593] &  i[1814]);
assign l_38[1818]    = ( l_39 [2594] & !i[1814]) | ( l_39 [2595] &  i[1814]);
assign l_38[1819]    = ( l_39 [2596] & !i[1814]) | ( l_39 [2597] &  i[1814]);
assign l_38[1820]    = ( l_39 [2598] & !i[1814]) | ( l_39 [2599] &  i[1814]);
assign l_38[1821]    = ( l_39 [2600] & !i[1814]) | ( l_39 [2601] &  i[1814]);
assign l_38[1822]    = ( l_39 [2602] & !i[1814]) | ( l_39 [2603] &  i[1814]);
assign l_38[1823]    = ( l_39 [2604] & !i[1814]) | ( l_39 [2605] &  i[1814]);
assign l_38[1824]    = ( l_39 [2606] & !i[1814]) | ( l_39 [2607] &  i[1814]);
assign l_38[1825]    = ( l_39 [2608] & !i[1814]) | ( l_39 [2609] &  i[1814]);
assign l_38[1826]    = ( l_39 [2610] & !i[1814]) | ( l_39 [2611] &  i[1814]);
assign l_38[1827]    = ( l_39 [2612] & !i[1814]) | ( l_39 [2613] &  i[1814]);
assign l_38[1828]    = ( l_39 [2614] & !i[1814]) | ( l_39 [2615] &  i[1814]);
assign l_38[1829]    = ( l_39 [2616] & !i[1814]) | ( l_39 [2617] &  i[1814]);
assign l_38[1830]    = ( l_39 [2618] & !i[1814]) | ( l_39 [2619] &  i[1814]);
assign l_38[1831]    = ( l_39 [2620] & !i[1814]) | ( l_39 [2621] &  i[1814]);
assign l_38[1832]    = ( l_39 [2622] & !i[1814]) | ( l_39 [2623] &  i[1814]);
assign l_38[1833]    = ( l_39 [2624] & !i[1814]) | ( l_39 [2625] &  i[1814]);
assign l_38[1834]    = ( l_39 [2626] & !i[1814]) | ( l_39 [2627] &  i[1814]);
assign l_38[1835]    = ( l_39 [2628] & !i[1814]) | ( l_39 [2629] &  i[1814]);
assign l_38[1836]    = ( l_39 [2630] & !i[1814]) | ( l_39 [2631] &  i[1814]);
assign l_38[1837]    = ( l_39 [2632] & !i[1814]) | ( l_39 [2633] &  i[1814]);
assign l_38[1838]    = ( l_39 [2634] & !i[1814]) | ( l_39 [2635] &  i[1814]);
assign l_38[1839]    = ( l_39 [2636] & !i[1814]) | ( l_39 [2637] &  i[1814]);
assign l_38[1840]    = ( l_39 [2638] & !i[1814]) | ( l_39 [2639] &  i[1814]);
assign l_38[1841]    = ( l_39 [2640] & !i[1814]) | ( l_39 [2641] &  i[1814]);
assign l_38[1842]    = ( l_39 [2642] & !i[1814]) | ( l_39 [2643] &  i[1814]);
assign l_38[1843]    = ( l_39 [2644] & !i[1814]) | ( l_39 [2645] &  i[1814]);
assign l_38[1844]    = ( l_39 [2646] & !i[1814]) | ( l_39 [2647] &  i[1814]);
assign l_38[1845]    = ( l_39 [2648] & !i[1814]) | ( l_39 [2649] &  i[1814]);
assign l_38[1846]    = ( l_39 [2650] & !i[1814]) | ( l_39 [2651] &  i[1814]);
assign l_38[1847]    = ( l_39 [2652] & !i[1814]) | ( l_39 [2653] &  i[1814]);
assign l_38[1848]    = ( l_39 [2654] & !i[1814]) | ( l_39 [2655] &  i[1814]);
assign l_38[1849]    = ( l_39 [2656] & !i[1814]) | ( l_39 [2657] &  i[1814]);
assign l_38[1850]    = ( l_39 [2658] & !i[1814]) | ( l_39 [2659] &  i[1814]);
assign l_38[1851]    = ( l_39 [2660] & !i[1814]) | ( l_39 [2661] &  i[1814]);
assign l_38[1852]    = ( l_39 [2662] & !i[1814]) | ( l_39 [2663] &  i[1814]);
assign l_38[1853]    = ( l_39 [2664] & !i[1814]) | ( l_39 [2665] &  i[1814]);
assign l_38[1854]    = ( l_39 [2666] & !i[1814]) | ( l_39 [2667] &  i[1814]);
assign l_38[1855]    = ( l_39 [2668] & !i[1814]) | ( l_39 [2669] &  i[1814]);
assign l_38[1856]    = ( l_39 [2670] & !i[1814]) | ( l_39 [2671] &  i[1814]);
assign l_38[1857]    = ( l_39 [2672] & !i[1814]) | ( l_39 [2673] &  i[1814]);
assign l_38[1858]    = ( l_39 [2674] & !i[1814]) | ( l_39 [2675] &  i[1814]);
assign l_38[1859]    = ( l_39 [2676] & !i[1814]) | ( l_39 [2677] &  i[1814]);
assign l_38[1860]    = ( l_39 [2678] & !i[1814]) | ( l_39 [2679] &  i[1814]);
assign l_38[1861]    = ( l_39 [2680] & !i[1814]) | ( l_39 [2681] &  i[1814]);
assign l_38[1862]    = ( l_39 [2682] & !i[1814]) | ( l_39 [2683] &  i[1814]);
assign l_38[1863]    = ( l_39 [2684] & !i[1814]) | ( l_39 [2685] &  i[1814]);
assign l_38[1864]    = ( l_39 [2686] & !i[1814]) | ( l_39 [2687] &  i[1814]);
assign l_38[1865]    = ( l_39 [2688] & !i[1814]) | ( l_39 [2689] &  i[1814]);
assign l_38[1866]    = ( l_39 [2690] & !i[1814]) | ( l_39 [2691] &  i[1814]);
assign l_38[1867]    = ( l_39 [2692] & !i[1814]) | ( l_39 [2693] &  i[1814]);
assign l_38[1868]    = ( l_39 [2694] & !i[1814]) | ( l_39 [2695] &  i[1814]);
assign l_38[1869]    = ( l_39 [2696] & !i[1814]) | ( l_39 [2697] &  i[1814]);
assign l_38[1870]    = ( l_39 [2698] & !i[1814]) | ( l_39 [2699] &  i[1814]);
assign l_38[1871]    = ( l_39 [2700] & !i[1814]) | ( l_39 [2701] &  i[1814]);
assign l_38[1872]    = ( l_39 [2702] & !i[1814]) | ( l_39 [2703] &  i[1814]);
assign l_38[1873]    = ( l_39 [2704] & !i[1814]) | ( l_39 [2705] &  i[1814]);
assign l_38[1874]    = ( l_39 [2706] & !i[1814]) | ( l_39 [2707] &  i[1814]);
assign l_38[1875]    = ( l_39 [2708] & !i[1814]) | ( l_39 [2709] &  i[1814]);
assign l_38[1876]    = ( l_39 [2710] & !i[1814]) | ( l_39 [2711] &  i[1814]);
assign l_38[1877]    = ( l_39 [2712] & !i[1814]) | ( l_39 [2713] &  i[1814]);
assign l_38[1878]    = ( l_39 [2714] & !i[1814]) | ( l_39 [2715] &  i[1814]);
assign l_38[1879]    = ( l_39 [2716] & !i[1814]) | ( l_39 [2717] &  i[1814]);
assign l_38[1880]    = ( l_39 [2718] & !i[1814]) | ( l_39 [2719] &  i[1814]);
assign l_38[1881]    = ( l_39 [2720] & !i[1814]) | ( l_39 [2721] &  i[1814]);
assign l_38[1882]    = ( l_39 [2722] & !i[1814]) | ( l_39 [2723] &  i[1814]);
assign l_38[1883]    = ( l_39 [2724] & !i[1814]) | ( l_39 [2725] &  i[1814]);
assign l_38[1884]    = ( l_39 [2726] & !i[1814]) | ( l_39 [2727] &  i[1814]);
assign l_38[1885]    = ( l_39 [2728] & !i[1814]) | ( l_39 [2729] &  i[1814]);
assign l_38[1886]    = ( l_39 [2730] & !i[1814]) | ( l_39 [2731] &  i[1814]);
assign l_38[1887]    = ( l_39 [2732] & !i[1814]) | ( l_39 [2733] &  i[1814]);
assign l_38[1888]    = ( l_39 [2734] & !i[1814]) | ( l_39 [2735] &  i[1814]);
assign l_38[1889]    = ( l_39 [2736] & !i[1814]) | ( l_39 [2737] &  i[1814]);
assign l_38[1890]    = ( l_39 [2738] & !i[1814]) | ( l_39 [2739] &  i[1814]);
assign l_38[1891]    = ( l_39 [2740] & !i[1814]) | ( l_39 [2741] &  i[1814]);
assign l_38[1892]    = ( l_39 [2742] & !i[1814]) | ( l_39 [2743] &  i[1814]);
assign l_38[1893]    = ( l_39 [2744] & !i[1814]) | ( l_39 [2745] &  i[1814]);
assign l_38[1894]    = ( l_39 [2746] & !i[1814]) | ( l_39 [2747] &  i[1814]);
assign l_38[1895]    = ( l_39 [2748] & !i[1814]) | ( l_39 [2749] &  i[1814]);
assign l_38[1896]    = ( l_39 [2750] & !i[1814]) | ( l_39 [2751] &  i[1814]);
assign l_38[1897]    = ( l_39 [2752] & !i[1814]) | ( l_39 [2753] &  i[1814]);
assign l_38[1898]    = ( l_39 [2754] & !i[1814]) | ( l_39 [2755] &  i[1814]);
assign l_38[1899]    = ( l_39 [2756] & !i[1814]) | ( l_39 [2757] &  i[1814]);
assign l_38[1900]    = ( l_39 [2758] & !i[1814]) | ( l_39 [2759] &  i[1814]);
assign l_38[1901]    = ( l_39 [2760] & !i[1814]) | ( l_39 [2761] &  i[1814]);
assign l_38[1902]    = ( l_39 [2762] & !i[1814]) | ( l_39 [2763] &  i[1814]);
assign l_38[1903]    = ( l_39 [2764] & !i[1814]) | ( l_39 [2765] &  i[1814]);
assign l_38[1904]    = ( l_39 [2766] & !i[1814]) | ( l_39 [2767] &  i[1814]);
assign l_38[1905]    = ( l_39 [2768] & !i[1814]) | ( l_39 [2769] &  i[1814]);
assign l_38[1906]    = ( l_39 [2770] & !i[1814]) | ( l_39 [2771] &  i[1814]);
assign l_38[1907]    = ( l_39 [2772] & !i[1814]) | ( l_39 [2773] &  i[1814]);
assign l_38[1908]    = ( l_39 [2774] & !i[1814]) | ( l_39 [2775] &  i[1814]);
assign l_38[1909]    = ( l_39 [2776] & !i[1814]) | ( l_39 [2777] &  i[1814]);
assign l_38[1910]    = ( l_39 [2778] & !i[1814]) | ( l_39 [2779] &  i[1814]);
assign l_38[1911]    = ( l_39 [2780] & !i[1814]) | ( l_39 [2781] &  i[1814]);
assign l_38[1912]    = ( l_39 [2782] & !i[1814]) | ( l_39 [2783] &  i[1814]);
assign l_38[1913]    = ( l_39 [2784] & !i[1814]) | ( l_39 [2785] &  i[1814]);
assign l_38[1914]    = ( l_39 [2786] & !i[1814]) | ( l_39 [2787] &  i[1814]);
assign l_38[1915]    = ( l_39 [2788] & !i[1814]) | ( l_39 [2789] &  i[1814]);
assign l_38[1916]    = ( l_39 [2790] & !i[1814]) | ( l_39 [2791] &  i[1814]);
assign l_38[1917]    = ( l_39 [2792] & !i[1814]) | ( l_39 [2793] &  i[1814]);
assign l_38[1918]    = ( l_39 [2794] & !i[1814]) | ( l_39 [2795] &  i[1814]);
assign l_38[1919]    = ( l_39 [2796] & !i[1814]) | ( l_39 [2797] &  i[1814]);
assign l_38[1920]    = ( l_39 [2798] & !i[1814]) | ( l_39 [2799] &  i[1814]);
assign l_38[1921]    = ( l_39 [2800] & !i[1814]) | ( l_39 [2801] &  i[1814]);
assign l_38[1922]    = ( l_39 [2802] & !i[1814]) | ( l_39 [2803] &  i[1814]);
assign l_38[1923]    = ( l_39 [2804] & !i[1814]) | ( l_39 [2805] &  i[1814]);
assign l_38[1924]    = ( l_39 [2806] & !i[1814]) | ( l_39 [2807] &  i[1814]);
assign l_38[1925]    = ( l_39 [2808] & !i[1814]) | ( l_39 [2809] &  i[1814]);
assign l_38[1926]    = ( l_39 [2810] & !i[1814]) | ( l_39 [2811] &  i[1814]);
assign l_38[1927]    = ( l_39 [2812] & !i[1814]) | ( l_39 [2813] &  i[1814]);
assign l_38[1928]    = ( l_39 [2814] & !i[1814]) | ( l_39 [2815] &  i[1814]);
assign l_38[1929]    = ( l_39 [2816] & !i[1814]) | ( l_39 [2817] &  i[1814]);
assign l_38[1930]    = ( l_39 [2818] & !i[1814]) | ( l_39 [2819] &  i[1814]);
assign l_38[1931]    = ( l_39 [2820] & !i[1814]) | ( l_39 [2821] &  i[1814]);
assign l_38[1932]    = ( l_39 [2822] & !i[1814]) | ( l_39 [2823] &  i[1814]);
assign l_38[1933]    = ( l_39 [2824] & !i[1814]) | ( l_39 [2825] &  i[1814]);
assign l_38[1934]    = ( l_39 [2826] & !i[1814]) | ( l_39 [2827] &  i[1814]);
assign l_38[1935]    = ( l_39 [2828] & !i[1814]) | ( l_39 [2829] &  i[1814]);
assign l_38[1936]    = ( l_39 [2830] & !i[1814]) | ( l_39 [2831] &  i[1814]);
assign l_38[1937]    = ( l_39 [2832] & !i[1814]) | ( l_39 [2833] &  i[1814]);
assign l_38[1938]    = ( l_39 [2834] & !i[1814]) | ( l_39 [2835] &  i[1814]);
assign l_38[1939]    = ( l_39 [2836] & !i[1814]) | ( l_39 [2837] &  i[1814]);
assign l_38[1940]    = ( l_39 [2838] & !i[1814]) | ( l_39 [2839] &  i[1814]);
assign l_38[1941]    = ( l_39 [2840] & !i[1814]) | ( l_39 [2841] &  i[1814]);
assign l_38[1942]    = ( l_39 [2842] & !i[1814]) | ( l_39 [2843] &  i[1814]);
assign l_38[1943]    = ( l_39 [2844] & !i[1814]) | ( l_39 [2845] &  i[1814]);
assign l_38[1944]    = ( l_39 [2846] & !i[1814]) | ( l_39 [2847] &  i[1814]);
assign l_38[1945]    = ( l_39 [2848] & !i[1814]) | ( l_39 [2849] &  i[1814]);
assign l_38[1946]    = ( l_39 [2850] & !i[1814]) | ( l_39 [2851] &  i[1814]);
assign l_38[1947]    = ( l_39 [2852] & !i[1814]) | ( l_39 [2853] &  i[1814]);
assign l_38[1948]    = ( l_39 [2854] & !i[1814]) | ( l_39 [2855] &  i[1814]);
assign l_38[1949]    = ( l_39 [2856] & !i[1814]) | ( l_39 [2857] &  i[1814]);
assign l_38[1950]    = ( l_39 [2858] & !i[1814]) | ( l_39 [2859] &  i[1814]);
assign l_38[1951]    = ( l_39 [2860] & !i[1814]) | ( l_39 [2861] &  i[1814]);
assign l_38[1952]    = ( l_39 [2862] & !i[1814]) | ( l_39 [2863] &  i[1814]);
assign l_38[1953]    = ( l_39 [2864] & !i[1814]) | ( l_39 [2865] &  i[1814]);
assign l_38[1954]    = ( l_39 [2866] & !i[1814]) | ( l_39 [2867] &  i[1814]);
assign l_38[1955]    = ( l_39 [2868] & !i[1814]) | ( l_39 [2869] &  i[1814]);
assign l_38[1956]    = ( l_39 [2870] & !i[1814]) | ( l_39 [2871] &  i[1814]);
assign l_38[1957]    = ( l_39 [2872] & !i[1814]) | ( l_39 [2873] &  i[1814]);
assign l_38[1958]    = ( l_39 [2874] & !i[1814]) | ( l_39 [2875] &  i[1814]);
assign l_38[1959]    = ( l_39 [2876] & !i[1814]) | ( l_39 [2877] &  i[1814]);
assign l_38[1960]    = ( l_39 [2878] & !i[1814]) | ( l_39 [2879] &  i[1814]);
assign l_38[1961]    = ( l_39 [2880] & !i[1814]) | ( l_39 [2881] &  i[1814]);
assign l_38[1962]    = ( l_39 [2882] & !i[1814]) | ( l_39 [2883] &  i[1814]);
assign l_38[1963]    = ( l_39 [2884] & !i[1814]) | ( l_39 [2885] &  i[1814]);
assign l_38[1964]    = ( l_39 [2886] & !i[1814]) | ( l_39 [2887] &  i[1814]);
assign l_38[1965]    = ( l_39 [2888] & !i[1814]) | ( l_39 [2889] &  i[1814]);
assign l_38[1966]    = ( l_39 [2890] & !i[1814]) | ( l_39 [2891] &  i[1814]);
assign l_38[1967]    = ( l_39 [2892] & !i[1814]) | ( l_39 [2893] &  i[1814]);
assign l_38[1968]    = ( l_39 [2894] & !i[1814]) | ( l_39 [2895] &  i[1814]);
assign l_38[1969]    = ( l_39 [2896] & !i[1814]) | ( l_39 [2897] &  i[1814]);
assign l_38[1970]    = ( l_39 [2898] & !i[1814]) | ( l_39 [2899] &  i[1814]);
assign l_38[1971]    = ( l_39 [2900] & !i[1814]) | ( l_39 [2901] &  i[1814]);
assign l_38[1972]    = ( l_39 [2902] & !i[1814]) | ( l_39 [2903] &  i[1814]);
assign l_38[1973]    = ( l_39 [2904] & !i[1814]) | ( l_39 [2905] &  i[1814]);
assign l_38[1974]    = ( l_39 [2906] & !i[1814]) | ( l_39 [2907] &  i[1814]);
assign l_38[1975]    = ( l_39 [2908] & !i[1814]) | ( l_39 [2909] &  i[1814]);
assign l_38[1976]    = ( l_39 [2910] & !i[1814]) | ( l_39 [2911] &  i[1814]);
assign l_38[1977]    = ( l_39 [2912] & !i[1814]) | ( l_39 [2913] &  i[1814]);
assign l_38[1978]    = ( l_39 [2914] & !i[1814]) | ( l_39 [2915] &  i[1814]);
assign l_38[1979]    = ( l_39 [2916] & !i[1814]) | ( l_39 [2917] &  i[1814]);
assign l_38[1980]    = ( l_39 [2918] & !i[1814]) | ( l_39 [2919] &  i[1814]);
assign l_38[1981]    = ( l_39 [2920] & !i[1814]) | ( l_39 [2921] &  i[1814]);
assign l_38[1982]    = ( l_39 [2922] & !i[1814]) | ( l_39 [2923] &  i[1814]);
assign l_38[1983]    = ( l_39 [2924] & !i[1814]) | ( l_39 [2925] &  i[1814]);
assign l_38[1984]    = ( l_39 [2926] & !i[1814]) | ( l_39 [2927] &  i[1814]);
assign l_38[1985]    = ( l_39 [2928] & !i[1814]) | ( l_39 [2929] &  i[1814]);
assign l_38[1986]    = ( l_39 [2930] & !i[1814]) | ( l_39 [2931] &  i[1814]);
assign l_38[1987]    = ( l_39 [2932] & !i[1814]) | ( l_39 [2933] &  i[1814]);
assign l_38[1988]    = ( l_39 [2934] & !i[1814]) | ( l_39 [2935] &  i[1814]);
assign l_38[1989]    = ( l_39 [2936] & !i[1814]) | ( l_39 [2937] &  i[1814]);
assign l_38[1990]    = ( l_39 [2938] & !i[1814]) | ( l_39 [2939] &  i[1814]);
assign l_38[1991]    = ( l_39 [2940] & !i[1814]) | ( l_39 [2941] &  i[1814]);
assign l_38[1992]    = ( l_39 [2942] & !i[1814]) | ( l_39 [2943] &  i[1814]);
assign l_38[1993]    = ( l_39 [2944] & !i[1814]) | ( l_39 [2945] &  i[1814]);
assign l_38[1994]    = ( l_39 [2946] & !i[1814]) | ( l_39 [2947] &  i[1814]);
assign l_38[1995]    = ( l_39 [2948] & !i[1814]) | ( l_39 [2949] &  i[1814]);
assign l_38[1996]    = ( l_39 [2950] & !i[1814]) | ( l_39 [2951] &  i[1814]);
assign l_38[1997]    = ( l_39 [2952] & !i[1814]) | ( l_39 [2953] &  i[1814]);
assign l_38[1998]    = ( l_39 [2954] & !i[1814]) | ( l_39 [2955] &  i[1814]);
assign l_38[1999]    = ( l_39 [2956] & !i[1814]) | ( l_39 [2957] &  i[1814]);
assign l_38[2000]    = ( l_39 [2958] & !i[1814]) | ( l_39 [2959] &  i[1814]);
assign l_38[2001]    = ( l_39 [2960] & !i[1814]) | ( l_39 [2961] &  i[1814]);
assign l_38[2002]    = ( l_39 [2962] & !i[1814]) | ( l_39 [2963] &  i[1814]);
assign l_38[2003]    = ( l_39 [2964] & !i[1814]) | ( l_39 [2965] &  i[1814]);
assign l_38[2004]    = ( l_39 [2966] & !i[1814]) | ( l_39 [2967] &  i[1814]);
assign l_38[2005]    = ( l_39 [2968] & !i[1814]) | ( l_39 [2969] &  i[1814]);
assign l_38[2006]    = ( l_39 [2970] & !i[1814]) | ( l_39 [2971] &  i[1814]);
assign l_38[2007]    = ( l_39 [2972] & !i[1814]) | ( l_39 [2973] &  i[1814]);
assign l_38[2008]    = ( l_39 [2974] & !i[1814]) | ( l_39 [2975] &  i[1814]);
assign l_38[2009]    = ( l_39 [2976] & !i[1814]) | ( l_39 [2977] &  i[1814]);
assign l_38[2010]    = ( l_39 [2978] & !i[1814]) | ( l_39 [2979] &  i[1814]);
assign l_38[2011]    = ( l_39 [2980] & !i[1814]) | ( l_39 [2981] &  i[1814]);
assign l_38[2012]    = ( l_39 [2982] & !i[1814]) | ( l_39 [2983] &  i[1814]);
assign l_38[2013]    = ( l_39 [2984] & !i[1814]) | ( l_39 [2985] &  i[1814]);
assign l_38[2014]    = ( l_39 [2986] & !i[1814]) | ( l_39 [2987] &  i[1814]);
assign l_38[2015]    = ( l_39 [2988] & !i[1814]) | ( l_39 [2989] &  i[1814]);
assign l_38[2016]    = ( l_39 [2990] & !i[1814]) | ( l_39 [2991] &  i[1814]);
assign l_38[2017]    = ( l_39 [2992] & !i[1814]) | ( l_39 [2993] &  i[1814]);
assign l_38[2018]    = ( l_39 [2994] & !i[1814]) | ( l_39 [2995] &  i[1814]);
assign l_38[2019]    = ( l_39 [2996] & !i[1814]) | ( l_39 [2997] &  i[1814]);
assign l_38[2020]    = ( l_39 [2998] & !i[1814]) | ( l_39 [2999] &  i[1814]);
assign l_38[2021]    = ( l_39 [3000] & !i[1814]) | ( l_39 [3001] &  i[1814]);
assign l_38[2022]    = ( l_39 [3002] & !i[1814]) | ( l_39 [3003] &  i[1814]);
assign l_38[2023]    = ( l_39 [3004] & !i[1814]) | ( l_39 [3005] &  i[1814]);
assign l_38[2024]    = ( l_39 [3006] & !i[1814]) | ( l_39 [3007] &  i[1814]);
assign l_38[2025]    = ( l_39 [3008] & !i[1814]) | ( l_39 [3009] &  i[1814]);
assign l_38[2026]    = ( l_39 [3010] & !i[1814]) | ( l_39 [3011] &  i[1814]);
assign l_38[2027]    = ( l_39 [3012] & !i[1814]) | ( l_39 [3013] &  i[1814]);
assign l_38[2028]    = ( l_39 [3014] & !i[1814]) | ( l_39 [3015] &  i[1814]);
assign l_38[2029]    = ( l_39 [3016] & !i[1814]) | ( l_39 [3017] &  i[1814]);
assign l_38[2030]    = ( l_39 [3018] & !i[1814]) | ( l_39 [3019] &  i[1814]);
assign l_38[2031]    = ( l_39 [3020] & !i[1814]) | ( l_39 [3021] &  i[1814]);
assign l_38[2032]    = ( l_39 [3022] & !i[1814]) | ( l_39 [3023] &  i[1814]);
assign l_38[2033]    = ( l_39 [3024] & !i[1814]) | ( l_39 [3025] &  i[1814]);
assign l_38[2034]    = ( l_39 [3026] & !i[1814]) | ( l_39 [3027] &  i[1814]);
assign l_38[2035]    = ( l_39 [3028] & !i[1814]) | ( l_39 [3029] &  i[1814]);
assign l_38[2036]    = ( l_39 [3030] & !i[1814]) | ( l_39 [3031] &  i[1814]);
assign l_38[2037]    = ( l_39 [3032] & !i[1814]) | ( l_39 [3033] &  i[1814]);
assign l_38[2038]    = ( l_39 [3034] & !i[1814]) | ( l_39 [3035] &  i[1814]);
assign l_38[2039]    = ( l_39 [3036] & !i[1814]) | ( l_39 [3037] &  i[1814]);
assign l_38[2040]    = ( l_39 [3038] & !i[1814]) | ( l_39 [3039] &  i[1814]);
assign l_38[2041]    = ( l_39 [3040] & !i[1814]) | ( l_39 [3041] &  i[1814]);
assign l_38[2042]    = ( l_39 [3042] & !i[1814]) | ( l_39 [3043] &  i[1814]);
assign l_38[2043]    = ( l_39 [3044] & !i[1814]) | ( l_39 [3045] &  i[1814]);
assign l_38[2044]    = ( l_39 [3046] & !i[1814]) | ( l_39 [3047] &  i[1814]);
assign l_38[2045]    = ( l_39 [3048] & !i[1814]) | ( l_39 [3049] &  i[1814]);
assign l_38[2046]    = ( l_39 [3050] & !i[1814]) | ( l_39 [3051] &  i[1814]);
assign l_38[2047]    = ( l_39 [3052] & !i[1814]) | ( l_39 [3053] &  i[1814]);
assign l_38[2048]    = ( l_39 [3054] & !i[1814]) | ( l_39 [3055] &  i[1814]);
assign l_38[2049]    = ( l_39 [3056] & !i[1814]) | ( l_39 [3057] &  i[1814]);
assign l_38[2050]    = ( l_39 [3058] & !i[1814]) | ( l_39 [3059] &  i[1814]);
assign l_38[2051]    = ( l_39 [3060] & !i[1814]) | ( l_39 [3061] &  i[1814]);
assign l_38[2052]    = ( l_39 [3062] & !i[1814]) | ( l_39 [3063] &  i[1814]);
assign l_38[2053]    = ( l_39 [3064] & !i[1814]) | ( l_39 [3065] &  i[1814]);
assign l_38[2054]    = ( l_39 [3066] & !i[1814]) | ( l_39 [3067] &  i[1814]);
assign l_38[2055]    = ( l_39 [3068] & !i[1814]) | ( l_39 [3069] &  i[1814]);
assign l_38[2056]    = ( l_39 [3070] & !i[1814]) | ( l_39 [3071] &  i[1814]);
assign l_38[2057]    = ( l_39 [3072] & !i[1814]) | ( l_39 [3073] &  i[1814]);
assign l_38[2058]    = ( l_39 [3074] & !i[1814]) | ( l_39 [3075] &  i[1814]);
assign l_38[2059]    = ( l_39 [3076] & !i[1814]) | ( l_39 [3077] &  i[1814]);
assign l_38[2060]    = ( l_39 [3078] & !i[1814]) | ( l_39 [3079] &  i[1814]);
assign l_38[2061]    = ( l_39 [3080] & !i[1814]) | ( l_39 [3081] &  i[1814]);
assign l_38[2062]    = ( l_39 [3082] & !i[1814]) | ( l_39 [3083] &  i[1814]);
assign l_38[2063]    = ( l_39 [3084] & !i[1814]) | ( l_39 [3085] &  i[1814]);
assign l_38[2064]    = ( l_39 [3086] & !i[1814]) | ( l_39 [3087] &  i[1814]);
assign l_38[2065]    = ( l_39 [3088] & !i[1814]) | ( l_39 [3089] &  i[1814]);
assign l_39[0]    = ( l_40 [0]);
assign l_39[1]    = ( l_40 [1] & !i[1817]);
assign l_39[2]    = ( l_40 [2] & !i[1817]);
assign l_39[3]    = (!i[1817]) | ( l_40 [3] &  i[1817]);
assign l_39[4]    = (!i[1817]) | ( l_40 [4] &  i[1817]);
assign l_39[5]    = ( l_40 [5] & !i[1817]);
assign l_39[6]    = ( l_40 [6] & !i[1817]);
assign l_39[7]    = (!i[1817]) | ( l_40 [7] &  i[1817]);
assign l_39[8]    = (!i[1817]) | ( l_40 [8] &  i[1817]);
assign l_39[9]    = ( l_40 [9] & !i[1817]) | ( l_40 [10] &  i[1817]);
assign l_39[10]    = ( l_40 [10]);
assign l_39[11]    = ( l_40 [11] & !i[1817]) | ( l_40 [10] &  i[1817]);
assign l_39[12]    = ( l_40 [10] & !i[1817]) | ( l_40 [12] &  i[1817]);
assign l_39[13]    = ( l_40 [10] & !i[1817]) | ( l_40 [13] &  i[1817]);
assign l_39[14]    = ( l_40 [14] & !i[1817]) | ( l_40 [10] &  i[1817]);
assign l_39[15]    = ( l_40 [15] & !i[1817]) | ( l_40 [10] &  i[1817]);
assign l_39[16]    = ( l_40 [10] & !i[1817]) | ( l_40 [16] &  i[1817]);
assign l_39[17]    = ( l_40 [10] & !i[1817]) | ( l_40 [17] &  i[1817]);
assign l_39[18]    = ( l_40 [18] & !i[1817]) | ( l_40 [19] &  i[1817]);
assign l_39[19]    = ( l_40 [20] & !i[1817]) | ( l_40 [21] &  i[1817]);
assign l_39[20]    = ( l_40 [22] & !i[1817]) | ( l_40 [23] &  i[1817]);
assign l_39[21]    = ( l_40 [24] & !i[1817]) | ( l_40 [25] &  i[1817]);
assign l_39[22]    = ( l_40 [26] & !i[1817]) | ( l_40 [27] &  i[1817]);
assign l_39[23]    = ( l_40 [28] & !i[1817]) | ( l_40 [29] &  i[1817]);
assign l_39[24]    = ( l_40 [30] & !i[1817]) | ( l_40 [31] &  i[1817]);
assign l_39[25]    = ( l_40 [32] & !i[1817]) | ( l_40 [33] &  i[1817]);
assign l_39[26]    = ( l_40 [34] & !i[1817]) | ( l_40 [35] &  i[1817]);
assign l_39[27]    = ( l_40 [36] & !i[1817]) | ( l_40 [37] &  i[1817]);
assign l_39[28]    = ( l_40 [38] & !i[1817]) | ( l_40 [39] &  i[1817]);
assign l_39[29]    = ( l_40 [40] & !i[1817]) | ( l_40 [41] &  i[1817]);
assign l_39[30]    = ( l_40 [42] & !i[1817]) | ( l_40 [43] &  i[1817]);
assign l_39[31]    = ( l_40 [44] & !i[1817]) | ( l_40 [45] &  i[1817]);
assign l_39[32]    = ( l_40 [46] & !i[1817]) | ( l_40 [47] &  i[1817]);
assign l_39[33]    = ( l_40 [48] & !i[1817]) | ( l_40 [49] &  i[1817]);
assign l_39[34]    = ( l_40 [50] & !i[1817]) | ( l_40 [51] &  i[1817]);
assign l_39[35]    = ( l_40 [52] & !i[1817]) | ( l_40 [53] &  i[1817]);
assign l_39[36]    = ( l_40 [54] & !i[1817]) | ( l_40 [55] &  i[1817]);
assign l_39[37]    = ( l_40 [56] & !i[1817]) | ( l_40 [57] &  i[1817]);
assign l_39[38]    = ( l_40 [58] & !i[1817]) | ( l_40 [59] &  i[1817]);
assign l_39[39]    = ( l_40 [60] & !i[1817]) | ( l_40 [61] &  i[1817]);
assign l_39[40]    = ( l_40 [62] & !i[1817]) | ( l_40 [63] &  i[1817]);
assign l_39[41]    = ( l_40 [64] & !i[1817]) | ( l_40 [65] &  i[1817]);
assign l_39[42]    = ( l_40 [66] & !i[1817]) | ( l_40 [67] &  i[1817]);
assign l_39[43]    = ( l_40 [68] & !i[1817]) | ( l_40 [69] &  i[1817]);
assign l_39[44]    = ( l_40 [70] & !i[1817]) | ( l_40 [71] &  i[1817]);
assign l_39[45]    = ( l_40 [72] & !i[1817]) | ( l_40 [73] &  i[1817]);
assign l_39[46]    = ( l_40 [74] & !i[1817]) | ( l_40 [75] &  i[1817]);
assign l_39[47]    = ( l_40 [76] & !i[1817]) | ( l_40 [77] &  i[1817]);
assign l_39[48]    = ( l_40 [78] & !i[1817]) | ( l_40 [79] &  i[1817]);
assign l_39[49]    = ( l_40 [80] & !i[1817]) | ( l_40 [81] &  i[1817]);
assign l_39[50]    = ( l_40 [82] & !i[1817]) | ( l_40 [83] &  i[1817]);
assign l_39[51]    = ( l_40 [84] & !i[1817]) | ( l_40 [85] &  i[1817]);
assign l_39[52]    = ( l_40 [86] & !i[1817]) | ( l_40 [87] &  i[1817]);
assign l_39[53]    = ( l_40 [88] & !i[1817]) | ( l_40 [89] &  i[1817]);
assign l_39[54]    = ( l_40 [90] & !i[1817]) | ( l_40 [91] &  i[1817]);
assign l_39[55]    = ( l_40 [92] & !i[1817]) | ( l_40 [93] &  i[1817]);
assign l_39[56]    = ( l_40 [94] & !i[1817]) | ( l_40 [95] &  i[1817]);
assign l_39[57]    = ( l_40 [96] & !i[1817]) | ( l_40 [97] &  i[1817]);
assign l_39[58]    = ( l_40 [98] & !i[1817]) | ( l_40 [99] &  i[1817]);
assign l_39[59]    = ( l_40 [100] & !i[1817]) | ( l_40 [101] &  i[1817]);
assign l_39[60]    = ( l_40 [102] & !i[1817]) | ( l_40 [103] &  i[1817]);
assign l_39[61]    = ( l_40 [104] & !i[1817]) | ( l_40 [105] &  i[1817]);
assign l_39[62]    = ( l_40 [106] & !i[1817]) | ( l_40 [107] &  i[1817]);
assign l_39[63]    = ( l_40 [108] & !i[1817]) | ( l_40 [109] &  i[1817]);
assign l_39[64]    = ( l_40 [110] & !i[1817]) | ( l_40 [111] &  i[1817]);
assign l_39[65]    = ( l_40 [112] & !i[1817]) | ( l_40 [113] &  i[1817]);
assign l_39[66]    = ( l_40 [114] & !i[1817]) | ( l_40 [115] &  i[1817]);
assign l_39[67]    = ( l_40 [116] & !i[1817]) | ( l_40 [117] &  i[1817]);
assign l_39[68]    = ( l_40 [118] & !i[1817]) | ( l_40 [119] &  i[1817]);
assign l_39[69]    = ( l_40 [120] & !i[1817]) | ( l_40 [121] &  i[1817]);
assign l_39[70]    = ( l_40 [122] & !i[1817]) | ( l_40 [123] &  i[1817]);
assign l_39[71]    = ( l_40 [124] & !i[1817]) | ( l_40 [125] &  i[1817]);
assign l_39[72]    = ( l_40 [126] & !i[1817]) | ( l_40 [127] &  i[1817]);
assign l_39[73]    = ( l_40 [128] & !i[1817]) | ( l_40 [129] &  i[1817]);
assign l_39[74]    = ( l_40 [130] & !i[1817]) | ( l_40 [131] &  i[1817]);
assign l_39[75]    = ( l_40 [132] & !i[1817]) | ( l_40 [133] &  i[1817]);
assign l_39[76]    = ( l_40 [134] & !i[1817]) | ( l_40 [135] &  i[1817]);
assign l_39[77]    = ( l_40 [136] & !i[1817]) | ( l_40 [137] &  i[1817]);
assign l_39[78]    = ( l_40 [138] & !i[1817]) | ( l_40 [139] &  i[1817]);
assign l_39[79]    = ( l_40 [140] & !i[1817]) | ( l_40 [141] &  i[1817]);
assign l_39[80]    = ( l_40 [142] & !i[1817]) | ( l_40 [143] &  i[1817]);
assign l_39[81]    = ( l_40 [144] & !i[1817]) | ( l_40 [145] &  i[1817]);
assign l_39[82]    = ( l_40 [146] & !i[1817]) | ( l_40 [147] &  i[1817]);
assign l_39[83]    = ( l_40 [148] & !i[1817]) | ( l_40 [149] &  i[1817]);
assign l_39[84]    = ( l_40 [150] & !i[1817]) | ( l_40 [151] &  i[1817]);
assign l_39[85]    = ( l_40 [152] & !i[1817]) | ( l_40 [153] &  i[1817]);
assign l_39[86]    = ( l_40 [154] & !i[1817]) | ( l_40 [155] &  i[1817]);
assign l_39[87]    = ( l_40 [156] & !i[1817]) | ( l_40 [157] &  i[1817]);
assign l_39[88]    = ( l_40 [158] & !i[1817]) | ( l_40 [159] &  i[1817]);
assign l_39[89]    = ( l_40 [160] & !i[1817]) | ( l_40 [161] &  i[1817]);
assign l_39[90]    = ( l_40 [162] & !i[1817]) | ( l_40 [163] &  i[1817]);
assign l_39[91]    = ( l_40 [164] & !i[1817]) | ( l_40 [165] &  i[1817]);
assign l_39[92]    = ( l_40 [166] & !i[1817]) | ( l_40 [167] &  i[1817]);
assign l_39[93]    = ( l_40 [168] & !i[1817]) | ( l_40 [169] &  i[1817]);
assign l_39[94]    = ( l_40 [170] & !i[1817]) | ( l_40 [171] &  i[1817]);
assign l_39[95]    = ( l_40 [172] & !i[1817]) | ( l_40 [173] &  i[1817]);
assign l_39[96]    = ( l_40 [174] & !i[1817]) | ( l_40 [175] &  i[1817]);
assign l_39[97]    = ( l_40 [176] & !i[1817]) | ( l_40 [177] &  i[1817]);
assign l_39[98]    = ( l_40 [178] & !i[1817]) | ( l_40 [179] &  i[1817]);
assign l_39[99]    = ( l_40 [180] & !i[1817]) | ( l_40 [181] &  i[1817]);
assign l_39[100]    = ( l_40 [182] & !i[1817]) | ( l_40 [183] &  i[1817]);
assign l_39[101]    = ( l_40 [184] & !i[1817]) | ( l_40 [185] &  i[1817]);
assign l_39[102]    = ( l_40 [186] & !i[1817]) | ( l_40 [187] &  i[1817]);
assign l_39[103]    = ( l_40 [188] & !i[1817]) | ( l_40 [189] &  i[1817]);
assign l_39[104]    = ( l_40 [190] & !i[1817]) | ( l_40 [191] &  i[1817]);
assign l_39[105]    = ( l_40 [192] & !i[1817]) | ( l_40 [193] &  i[1817]);
assign l_39[106]    = ( l_40 [194] & !i[1817]) | ( l_40 [195] &  i[1817]);
assign l_39[107]    = ( l_40 [196] & !i[1817]) | ( l_40 [197] &  i[1817]);
assign l_39[108]    = ( l_40 [198] & !i[1817]) | ( l_40 [199] &  i[1817]);
assign l_39[109]    = ( l_40 [200] & !i[1817]) | ( l_40 [201] &  i[1817]);
assign l_39[110]    = ( l_40 [202] & !i[1817]) | ( l_40 [203] &  i[1817]);
assign l_39[111]    = ( l_40 [204] & !i[1817]) | ( l_40 [205] &  i[1817]);
assign l_39[112]    = ( l_40 [206] & !i[1817]) | ( l_40 [207] &  i[1817]);
assign l_39[113]    = ( l_40 [208] & !i[1817]) | ( l_40 [209] &  i[1817]);
assign l_39[114]    = ( l_40 [210] & !i[1817]) | ( l_40 [211] &  i[1817]);
assign l_39[115]    = ( l_40 [212] & !i[1817]) | ( l_40 [213] &  i[1817]);
assign l_39[116]    = ( l_40 [214] & !i[1817]) | ( l_40 [215] &  i[1817]);
assign l_39[117]    = ( l_40 [216] & !i[1817]) | ( l_40 [217] &  i[1817]);
assign l_39[118]    = ( l_40 [218] & !i[1817]) | ( l_40 [219] &  i[1817]);
assign l_39[119]    = ( l_40 [220] & !i[1817]) | ( l_40 [221] &  i[1817]);
assign l_39[120]    = ( l_40 [222] & !i[1817]) | ( l_40 [223] &  i[1817]);
assign l_39[121]    = ( l_40 [224] & !i[1817]) | ( l_40 [225] &  i[1817]);
assign l_39[122]    = ( l_40 [226] & !i[1817]) | ( l_40 [227] &  i[1817]);
assign l_39[123]    = ( l_40 [228] & !i[1817]) | ( l_40 [229] &  i[1817]);
assign l_39[124]    = ( l_40 [230] & !i[1817]) | ( l_40 [231] &  i[1817]);
assign l_39[125]    = ( l_40 [232] & !i[1817]) | ( l_40 [233] &  i[1817]);
assign l_39[126]    = ( l_40 [234] & !i[1817]) | ( l_40 [235] &  i[1817]);
assign l_39[127]    = ( l_40 [236] & !i[1817]) | ( l_40 [237] &  i[1817]);
assign l_39[128]    = ( l_40 [238] & !i[1817]) | ( l_40 [239] &  i[1817]);
assign l_39[129]    = ( l_40 [240] & !i[1817]) | ( l_40 [241] &  i[1817]);
assign l_39[130]    = ( l_40 [242] & !i[1817]) | ( l_40 [243] &  i[1817]);
assign l_39[131]    = ( l_40 [244] & !i[1817]) | ( l_40 [245] &  i[1817]);
assign l_39[132]    = ( l_40 [246] & !i[1817]) | ( l_40 [247] &  i[1817]);
assign l_39[133]    = ( l_40 [248] & !i[1817]) | ( l_40 [249] &  i[1817]);
assign l_39[134]    = ( l_40 [250] & !i[1817]) | ( l_40 [251] &  i[1817]);
assign l_39[135]    = ( l_40 [252] & !i[1817]) | ( l_40 [253] &  i[1817]);
assign l_39[136]    = ( l_40 [254] & !i[1817]) | ( l_40 [255] &  i[1817]);
assign l_39[137]    = ( l_40 [256] & !i[1817]) | ( l_40 [257] &  i[1817]);
assign l_39[138]    = ( l_40 [258] & !i[1817]) | ( l_40 [259] &  i[1817]);
assign l_39[139]    = ( l_40 [260] & !i[1817]) | ( l_40 [261] &  i[1817]);
assign l_39[140]    = ( l_40 [262] & !i[1817]) | ( l_40 [263] &  i[1817]);
assign l_39[141]    = ( l_40 [264] & !i[1817]) | ( l_40 [265] &  i[1817]);
assign l_39[142]    = ( l_40 [266] & !i[1817]) | ( l_40 [267] &  i[1817]);
assign l_39[143]    = ( l_40 [268] & !i[1817]) | ( l_40 [269] &  i[1817]);
assign l_39[144]    = ( l_40 [270] & !i[1817]) | ( l_40 [271] &  i[1817]);
assign l_39[145]    = ( l_40 [272] & !i[1817]) | ( l_40 [273] &  i[1817]);
assign l_39[146]    = ( l_40 [274] & !i[1817]) | ( l_40 [275] &  i[1817]);
assign l_39[147]    = ( l_40 [276] & !i[1817]) | ( l_40 [277] &  i[1817]);
assign l_39[148]    = ( l_40 [278] & !i[1817]) | ( l_40 [279] &  i[1817]);
assign l_39[149]    = ( l_40 [280] & !i[1817]) | ( l_40 [281] &  i[1817]);
assign l_39[150]    = ( l_40 [282] & !i[1817]) | ( l_40 [283] &  i[1817]);
assign l_39[151]    = ( l_40 [284] & !i[1817]) | ( l_40 [285] &  i[1817]);
assign l_39[152]    = ( l_40 [286] & !i[1817]) | ( l_40 [287] &  i[1817]);
assign l_39[153]    = ( l_40 [288] & !i[1817]) | ( l_40 [289] &  i[1817]);
assign l_39[154]    = ( l_40 [290] & !i[1817]) | ( l_40 [291] &  i[1817]);
assign l_39[155]    = ( l_40 [292] & !i[1817]) | ( l_40 [293] &  i[1817]);
assign l_39[156]    = ( l_40 [294] & !i[1817]) | ( l_40 [295] &  i[1817]);
assign l_39[157]    = ( l_40 [296] & !i[1817]) | ( l_40 [297] &  i[1817]);
assign l_39[158]    = ( l_40 [298] & !i[1817]) | ( l_40 [299] &  i[1817]);
assign l_39[159]    = ( l_40 [300] & !i[1817]) | ( l_40 [301] &  i[1817]);
assign l_39[160]    = ( l_40 [302] & !i[1817]) | ( l_40 [303] &  i[1817]);
assign l_39[161]    = ( l_40 [304] & !i[1817]) | ( l_40 [305] &  i[1817]);
assign l_39[162]    = ( l_40 [306] & !i[1817]) | ( l_40 [307] &  i[1817]);
assign l_39[163]    = ( l_40 [308] & !i[1817]) | ( l_40 [309] &  i[1817]);
assign l_39[164]    = ( l_40 [310] & !i[1817]) | ( l_40 [311] &  i[1817]);
assign l_39[165]    = ( l_40 [312] & !i[1817]) | ( l_40 [313] &  i[1817]);
assign l_39[166]    = ( l_40 [314] & !i[1817]) | ( l_40 [315] &  i[1817]);
assign l_39[167]    = ( l_40 [316] & !i[1817]) | ( l_40 [317] &  i[1817]);
assign l_39[168]    = ( l_40 [318] & !i[1817]) | ( l_40 [319] &  i[1817]);
assign l_39[169]    = ( l_40 [320] & !i[1817]) | ( l_40 [321] &  i[1817]);
assign l_39[170]    = ( l_40 [322] & !i[1817]) | ( l_40 [323] &  i[1817]);
assign l_39[171]    = ( l_40 [324] & !i[1817]) | ( l_40 [325] &  i[1817]);
assign l_39[172]    = ( l_40 [326] & !i[1817]) | ( l_40 [327] &  i[1817]);
assign l_39[173]    = ( l_40 [328] & !i[1817]) | ( l_40 [329] &  i[1817]);
assign l_39[174]    = ( l_40 [330] & !i[1817]) | ( l_40 [331] &  i[1817]);
assign l_39[175]    = ( l_40 [332] & !i[1817]) | ( l_40 [333] &  i[1817]);
assign l_39[176]    = ( l_40 [334] & !i[1817]) | ( l_40 [335] &  i[1817]);
assign l_39[177]    = ( l_40 [336] & !i[1817]) | ( l_40 [337] &  i[1817]);
assign l_39[178]    = ( l_40 [338] & !i[1817]) | ( l_40 [339] &  i[1817]);
assign l_39[179]    = ( l_40 [340] & !i[1817]) | ( l_40 [341] &  i[1817]);
assign l_39[180]    = ( l_40 [342] & !i[1817]) | ( l_40 [343] &  i[1817]);
assign l_39[181]    = ( l_40 [344] & !i[1817]) | ( l_40 [345] &  i[1817]);
assign l_39[182]    = ( l_40 [346] & !i[1817]) | ( l_40 [347] &  i[1817]);
assign l_39[183]    = ( l_40 [348] & !i[1817]) | ( l_40 [349] &  i[1817]);
assign l_39[184]    = ( l_40 [350] & !i[1817]) | ( l_40 [351] &  i[1817]);
assign l_39[185]    = ( l_40 [352] & !i[1817]) | ( l_40 [353] &  i[1817]);
assign l_39[186]    = ( l_40 [354] & !i[1817]) | ( l_40 [355] &  i[1817]);
assign l_39[187]    = ( l_40 [356] & !i[1817]) | ( l_40 [357] &  i[1817]);
assign l_39[188]    = ( l_40 [358] & !i[1817]) | ( l_40 [359] &  i[1817]);
assign l_39[189]    = ( l_40 [360] & !i[1817]) | ( l_40 [361] &  i[1817]);
assign l_39[190]    = ( l_40 [362] & !i[1817]) | ( l_40 [363] &  i[1817]);
assign l_39[191]    = ( l_40 [364] & !i[1817]) | ( l_40 [365] &  i[1817]);
assign l_39[192]    = ( l_40 [366] & !i[1817]) | ( l_40 [367] &  i[1817]);
assign l_39[193]    = ( l_40 [368] & !i[1817]) | ( l_40 [369] &  i[1817]);
assign l_39[194]    = ( l_40 [370] & !i[1817]) | ( l_40 [371] &  i[1817]);
assign l_39[195]    = ( l_40 [372] & !i[1817]) | ( l_40 [373] &  i[1817]);
assign l_39[196]    = ( l_40 [374] & !i[1817]) | ( l_40 [375] &  i[1817]);
assign l_39[197]    = ( l_40 [376] & !i[1817]) | ( l_40 [377] &  i[1817]);
assign l_39[198]    = ( l_40 [378] & !i[1817]) | ( l_40 [379] &  i[1817]);
assign l_39[199]    = ( l_40 [380] & !i[1817]) | ( l_40 [381] &  i[1817]);
assign l_39[200]    = ( l_40 [382] & !i[1817]) | ( l_40 [383] &  i[1817]);
assign l_39[201]    = ( l_40 [384] & !i[1817]) | ( l_40 [385] &  i[1817]);
assign l_39[202]    = ( l_40 [386] & !i[1817]) | ( l_40 [387] &  i[1817]);
assign l_39[203]    = ( l_40 [388] & !i[1817]) | ( l_40 [389] &  i[1817]);
assign l_39[204]    = ( l_40 [390] & !i[1817]) | ( l_40 [391] &  i[1817]);
assign l_39[205]    = ( l_40 [392] & !i[1817]) | ( l_40 [393] &  i[1817]);
assign l_39[206]    = ( l_40 [394] & !i[1817]) | ( l_40 [395] &  i[1817]);
assign l_39[207]    = ( l_40 [396] & !i[1817]) | ( l_40 [397] &  i[1817]);
assign l_39[208]    = ( l_40 [398] & !i[1817]) | ( l_40 [399] &  i[1817]);
assign l_39[209]    = ( l_40 [400] & !i[1817]) | ( l_40 [401] &  i[1817]);
assign l_39[210]    = ( l_40 [402] & !i[1817]) | ( l_40 [403] &  i[1817]);
assign l_39[211]    = ( l_40 [404] & !i[1817]) | ( l_40 [405] &  i[1817]);
assign l_39[212]    = ( l_40 [406] & !i[1817]) | ( l_40 [407] &  i[1817]);
assign l_39[213]    = ( l_40 [408] & !i[1817]) | ( l_40 [409] &  i[1817]);
assign l_39[214]    = ( l_40 [410] & !i[1817]) | ( l_40 [411] &  i[1817]);
assign l_39[215]    = ( l_40 [412] & !i[1817]) | ( l_40 [413] &  i[1817]);
assign l_39[216]    = ( l_40 [414] & !i[1817]) | ( l_40 [415] &  i[1817]);
assign l_39[217]    = ( l_40 [416] & !i[1817]) | ( l_40 [417] &  i[1817]);
assign l_39[218]    = ( l_40 [418] & !i[1817]) | ( l_40 [419] &  i[1817]);
assign l_39[219]    = ( l_40 [420] & !i[1817]) | ( l_40 [421] &  i[1817]);
assign l_39[220]    = ( l_40 [422] & !i[1817]) | ( l_40 [423] &  i[1817]);
assign l_39[221]    = ( l_40 [424] & !i[1817]) | ( l_40 [425] &  i[1817]);
assign l_39[222]    = ( l_40 [426] & !i[1817]) | ( l_40 [427] &  i[1817]);
assign l_39[223]    = ( l_40 [428] & !i[1817]) | ( l_40 [429] &  i[1817]);
assign l_39[224]    = ( l_40 [430] & !i[1817]) | ( l_40 [431] &  i[1817]);
assign l_39[225]    = ( l_40 [432] & !i[1817]) | ( l_40 [433] &  i[1817]);
assign l_39[226]    = ( l_40 [434] & !i[1817]) | ( l_40 [435] &  i[1817]);
assign l_39[227]    = ( l_40 [436] & !i[1817]) | ( l_40 [437] &  i[1817]);
assign l_39[228]    = ( l_40 [438] & !i[1817]) | ( l_40 [439] &  i[1817]);
assign l_39[229]    = ( l_40 [440] & !i[1817]) | ( l_40 [441] &  i[1817]);
assign l_39[230]    = ( l_40 [442] & !i[1817]) | ( l_40 [443] &  i[1817]);
assign l_39[231]    = ( l_40 [444] & !i[1817]) | ( l_40 [445] &  i[1817]);
assign l_39[232]    = ( l_40 [446] & !i[1817]) | ( l_40 [447] &  i[1817]);
assign l_39[233]    = ( l_40 [448] & !i[1817]) | ( l_40 [449] &  i[1817]);
assign l_39[234]    = ( l_40 [450] & !i[1817]) | ( l_40 [451] &  i[1817]);
assign l_39[235]    = ( l_40 [452] & !i[1817]) | ( l_40 [453] &  i[1817]);
assign l_39[236]    = ( l_40 [454] & !i[1817]) | ( l_40 [455] &  i[1817]);
assign l_39[237]    = ( l_40 [456] & !i[1817]) | ( l_40 [457] &  i[1817]);
assign l_39[238]    = ( l_40 [458] & !i[1817]) | ( l_40 [459] &  i[1817]);
assign l_39[239]    = ( l_40 [460] & !i[1817]) | ( l_40 [461] &  i[1817]);
assign l_39[240]    = ( l_40 [462] & !i[1817]) | ( l_40 [463] &  i[1817]);
assign l_39[241]    = ( l_40 [464] & !i[1817]) | ( l_40 [465] &  i[1817]);
assign l_39[242]    = ( l_40 [466] & !i[1817]) | ( l_40 [467] &  i[1817]);
assign l_39[243]    = ( l_40 [468] & !i[1817]) | ( l_40 [469] &  i[1817]);
assign l_39[244]    = ( l_40 [470] & !i[1817]) | ( l_40 [471] &  i[1817]);
assign l_39[245]    = ( l_40 [472] & !i[1817]) | ( l_40 [473] &  i[1817]);
assign l_39[246]    = ( l_40 [474] & !i[1817]) | ( l_40 [475] &  i[1817]);
assign l_39[247]    = ( l_40 [476] & !i[1817]) | ( l_40 [477] &  i[1817]);
assign l_39[248]    = ( l_40 [478] & !i[1817]) | ( l_40 [479] &  i[1817]);
assign l_39[249]    = ( l_40 [480] & !i[1817]) | ( l_40 [481] &  i[1817]);
assign l_39[250]    = ( l_40 [482] & !i[1817]) | ( l_40 [483] &  i[1817]);
assign l_39[251]    = ( l_40 [484] & !i[1817]) | ( l_40 [485] &  i[1817]);
assign l_39[252]    = ( l_40 [486] & !i[1817]) | ( l_40 [487] &  i[1817]);
assign l_39[253]    = ( l_40 [488] & !i[1817]) | ( l_40 [489] &  i[1817]);
assign l_39[254]    = ( l_40 [490] & !i[1817]) | ( l_40 [491] &  i[1817]);
assign l_39[255]    = ( l_40 [492] & !i[1817]) | ( l_40 [493] &  i[1817]);
assign l_39[256]    = ( l_40 [494] & !i[1817]) | ( l_40 [495] &  i[1817]);
assign l_39[257]    = ( l_40 [496] & !i[1817]) | ( l_40 [497] &  i[1817]);
assign l_39[258]    = ( l_40 [498] & !i[1817]) | ( l_40 [499] &  i[1817]);
assign l_39[259]    = ( l_40 [500] & !i[1817]) | ( l_40 [501] &  i[1817]);
assign l_39[260]    = ( l_40 [502] & !i[1817]) | ( l_40 [503] &  i[1817]);
assign l_39[261]    = ( l_40 [504] & !i[1817]) | ( l_40 [505] &  i[1817]);
assign l_39[262]    = ( l_40 [506] & !i[1817]) | ( l_40 [507] &  i[1817]);
assign l_39[263]    = ( l_40 [508] & !i[1817]) | ( l_40 [509] &  i[1817]);
assign l_39[264]    = ( l_40 [510] & !i[1817]) | ( l_40 [511] &  i[1817]);
assign l_39[265]    = ( l_40 [512] & !i[1817]) | ( l_40 [513] &  i[1817]);
assign l_39[266]    = ( l_40 [514] & !i[1817]) | ( l_40 [515] &  i[1817]);
assign l_39[267]    = ( l_40 [516] & !i[1817]) | ( l_40 [517] &  i[1817]);
assign l_39[268]    = ( l_40 [518] & !i[1817]) | ( l_40 [519] &  i[1817]);
assign l_39[269]    = ( l_40 [520] & !i[1817]) | ( l_40 [521] &  i[1817]);
assign l_39[270]    = ( l_40 [522] & !i[1817]) | ( l_40 [523] &  i[1817]);
assign l_39[271]    = ( l_40 [524] & !i[1817]) | ( l_40 [525] &  i[1817]);
assign l_39[272]    = ( l_40 [526] & !i[1817]) | ( l_40 [527] &  i[1817]);
assign l_39[273]    = ( l_40 [528] & !i[1817]) | ( l_40 [529] &  i[1817]);
assign l_39[274]    = ( l_40 [530] & !i[1817]) | ( l_40 [531] &  i[1817]);
assign l_39[275]    = ( l_40 [532] & !i[1817]) | ( l_40 [533] &  i[1817]);
assign l_39[276]    = ( l_40 [534] & !i[1817]) | ( l_40 [535] &  i[1817]);
assign l_39[277]    = ( l_40 [536] & !i[1817]) | ( l_40 [537] &  i[1817]);
assign l_39[278]    = ( l_40 [538] & !i[1817]) | ( l_40 [539] &  i[1817]);
assign l_39[279]    = ( l_40 [540] & !i[1817]) | ( l_40 [541] &  i[1817]);
assign l_39[280]    = ( l_40 [542] & !i[1817]) | ( l_40 [543] &  i[1817]);
assign l_39[281]    = ( l_40 [544] & !i[1817]) | ( l_40 [545] &  i[1817]);
assign l_39[282]    = ( l_40 [546] & !i[1817]) | ( l_40 [547] &  i[1817]);
assign l_39[283]    = ( l_40 [548] & !i[1817]) | ( l_40 [549] &  i[1817]);
assign l_39[284]    = ( l_40 [550] & !i[1817]) | ( l_40 [551] &  i[1817]);
assign l_39[285]    = ( l_40 [552] & !i[1817]) | ( l_40 [553] &  i[1817]);
assign l_39[286]    = ( l_40 [554] & !i[1817]) | ( l_40 [555] &  i[1817]);
assign l_39[287]    = ( l_40 [556] & !i[1817]) | ( l_40 [557] &  i[1817]);
assign l_39[288]    = ( l_40 [558] & !i[1817]) | ( l_40 [559] &  i[1817]);
assign l_39[289]    = ( l_40 [560] & !i[1817]) | ( l_40 [561] &  i[1817]);
assign l_39[290]    = ( l_40 [562] & !i[1817]) | ( l_40 [563] &  i[1817]);
assign l_39[291]    = ( l_40 [564] & !i[1817]) | ( l_40 [565] &  i[1817]);
assign l_39[292]    = ( l_40 [566] & !i[1817]) | ( l_40 [567] &  i[1817]);
assign l_39[293]    = ( l_40 [568] & !i[1817]) | ( l_40 [569] &  i[1817]);
assign l_39[294]    = ( l_40 [570] & !i[1817]) | ( l_40 [571] &  i[1817]);
assign l_39[295]    = ( l_40 [572] & !i[1817]) | ( l_40 [573] &  i[1817]);
assign l_39[296]    = ( l_40 [574] & !i[1817]) | ( l_40 [575] &  i[1817]);
assign l_39[297]    = ( l_40 [576] & !i[1817]) | ( l_40 [577] &  i[1817]);
assign l_39[298]    = ( l_40 [578] & !i[1817]) | ( l_40 [579] &  i[1817]);
assign l_39[299]    = ( l_40 [580] & !i[1817]) | ( l_40 [581] &  i[1817]);
assign l_39[300]    = ( l_40 [582] & !i[1817]) | ( l_40 [583] &  i[1817]);
assign l_39[301]    = ( l_40 [584] & !i[1817]) | ( l_40 [585] &  i[1817]);
assign l_39[302]    = ( l_40 [586] & !i[1817]) | ( l_40 [587] &  i[1817]);
assign l_39[303]    = ( l_40 [588] & !i[1817]) | ( l_40 [589] &  i[1817]);
assign l_39[304]    = ( l_40 [590] & !i[1817]) | ( l_40 [591] &  i[1817]);
assign l_39[305]    = ( l_40 [592] & !i[1817]) | ( l_40 [593] &  i[1817]);
assign l_39[306]    = ( l_40 [594] & !i[1817]) | ( l_40 [595] &  i[1817]);
assign l_39[307]    = ( l_40 [596] & !i[1817]) | ( l_40 [597] &  i[1817]);
assign l_39[308]    = ( l_40 [598] & !i[1817]) | ( l_40 [599] &  i[1817]);
assign l_39[309]    = ( l_40 [600] & !i[1817]) | ( l_40 [601] &  i[1817]);
assign l_39[310]    = ( l_40 [602] & !i[1817]) | ( l_40 [603] &  i[1817]);
assign l_39[311]    = ( l_40 [604] & !i[1817]) | ( l_40 [605] &  i[1817]);
assign l_39[312]    = ( l_40 [606] & !i[1817]) | ( l_40 [607] &  i[1817]);
assign l_39[313]    = ( l_40 [608] & !i[1817]) | ( l_40 [609] &  i[1817]);
assign l_39[314]    = ( l_40 [610] & !i[1817]) | ( l_40 [611] &  i[1817]);
assign l_39[315]    = ( l_40 [612] & !i[1817]) | ( l_40 [613] &  i[1817]);
assign l_39[316]    = ( l_40 [614] & !i[1817]) | ( l_40 [615] &  i[1817]);
assign l_39[317]    = ( l_40 [616] & !i[1817]) | ( l_40 [617] &  i[1817]);
assign l_39[318]    = ( l_40 [618] & !i[1817]) | ( l_40 [619] &  i[1817]);
assign l_39[319]    = ( l_40 [620] & !i[1817]) | ( l_40 [621] &  i[1817]);
assign l_39[320]    = ( l_40 [622] & !i[1817]) | ( l_40 [623] &  i[1817]);
assign l_39[321]    = ( l_40 [624] & !i[1817]) | ( l_40 [625] &  i[1817]);
assign l_39[322]    = ( l_40 [626] & !i[1817]) | ( l_40 [627] &  i[1817]);
assign l_39[323]    = ( l_40 [628] & !i[1817]) | ( l_40 [629] &  i[1817]);
assign l_39[324]    = ( l_40 [630] & !i[1817]) | ( l_40 [631] &  i[1817]);
assign l_39[325]    = ( l_40 [632] & !i[1817]) | ( l_40 [633] &  i[1817]);
assign l_39[326]    = ( l_40 [634] & !i[1817]) | ( l_40 [635] &  i[1817]);
assign l_39[327]    = ( l_40 [636] & !i[1817]) | ( l_40 [637] &  i[1817]);
assign l_39[328]    = ( l_40 [638] & !i[1817]) | ( l_40 [639] &  i[1817]);
assign l_39[329]    = ( l_40 [640] & !i[1817]) | ( l_40 [641] &  i[1817]);
assign l_39[330]    = ( l_40 [642] & !i[1817]) | ( l_40 [643] &  i[1817]);
assign l_39[331]    = ( l_40 [644] & !i[1817]) | ( l_40 [645] &  i[1817]);
assign l_39[332]    = ( l_40 [646] & !i[1817]) | ( l_40 [647] &  i[1817]);
assign l_39[333]    = ( l_40 [648] & !i[1817]) | ( l_40 [649] &  i[1817]);
assign l_39[334]    = ( l_40 [650] & !i[1817]) | ( l_40 [651] &  i[1817]);
assign l_39[335]    = ( l_40 [652] & !i[1817]) | ( l_40 [653] &  i[1817]);
assign l_39[336]    = ( l_40 [654] & !i[1817]) | ( l_40 [655] &  i[1817]);
assign l_39[337]    = ( l_40 [656] & !i[1817]) | ( l_40 [657] &  i[1817]);
assign l_39[338]    = ( l_40 [658] & !i[1817]) | ( l_40 [659] &  i[1817]);
assign l_39[339]    = ( l_40 [660] & !i[1817]) | ( l_40 [661] &  i[1817]);
assign l_39[340]    = ( l_40 [662] & !i[1817]) | ( l_40 [663] &  i[1817]);
assign l_39[341]    = ( l_40 [664] & !i[1817]) | ( l_40 [665] &  i[1817]);
assign l_39[342]    = ( l_40 [666] & !i[1817]) | ( l_40 [667] &  i[1817]);
assign l_39[343]    = ( l_40 [668] & !i[1817]) | ( l_40 [669] &  i[1817]);
assign l_39[344]    = ( l_40 [670] & !i[1817]) | ( l_40 [671] &  i[1817]);
assign l_39[345]    = ( l_40 [672] & !i[1817]) | ( l_40 [673] &  i[1817]);
assign l_39[346]    = ( l_40 [674] & !i[1817]) | ( l_40 [675] &  i[1817]);
assign l_39[347]    = ( l_40 [676] & !i[1817]) | ( l_40 [677] &  i[1817]);
assign l_39[348]    = ( l_40 [678] & !i[1817]) | ( l_40 [679] &  i[1817]);
assign l_39[349]    = ( l_40 [680] & !i[1817]) | ( l_40 [681] &  i[1817]);
assign l_39[350]    = ( l_40 [682] & !i[1817]) | ( l_40 [683] &  i[1817]);
assign l_39[351]    = ( l_40 [684] & !i[1817]) | ( l_40 [685] &  i[1817]);
assign l_39[352]    = ( l_40 [686] & !i[1817]) | ( l_40 [687] &  i[1817]);
assign l_39[353]    = ( l_40 [688] & !i[1817]) | ( l_40 [689] &  i[1817]);
assign l_39[354]    = ( l_40 [690] & !i[1817]) | ( l_40 [691] &  i[1817]);
assign l_39[355]    = ( l_40 [692] & !i[1817]) | ( l_40 [693] &  i[1817]);
assign l_39[356]    = ( l_40 [694] & !i[1817]) | ( l_40 [695] &  i[1817]);
assign l_39[357]    = ( l_40 [696] & !i[1817]) | ( l_40 [697] &  i[1817]);
assign l_39[358]    = ( l_40 [698] & !i[1817]) | ( l_40 [699] &  i[1817]);
assign l_39[359]    = ( l_40 [700] & !i[1817]) | ( l_40 [701] &  i[1817]);
assign l_39[360]    = ( l_40 [702] & !i[1817]) | ( l_40 [703] &  i[1817]);
assign l_39[361]    = ( l_40 [704] & !i[1817]) | ( l_40 [705] &  i[1817]);
assign l_39[362]    = ( l_40 [706] & !i[1817]) | ( l_40 [707] &  i[1817]);
assign l_39[363]    = ( l_40 [708] & !i[1817]) | ( l_40 [709] &  i[1817]);
assign l_39[364]    = ( l_40 [710] & !i[1817]) | ( l_40 [711] &  i[1817]);
assign l_39[365]    = ( l_40 [712] & !i[1817]) | ( l_40 [713] &  i[1817]);
assign l_39[366]    = ( l_40 [714] & !i[1817]) | ( l_40 [715] &  i[1817]);
assign l_39[367]    = ( l_40 [716] & !i[1817]) | ( l_40 [717] &  i[1817]);
assign l_39[368]    = ( l_40 [718] & !i[1817]) | ( l_40 [719] &  i[1817]);
assign l_39[369]    = ( l_40 [720] & !i[1817]) | ( l_40 [721] &  i[1817]);
assign l_39[370]    = ( l_40 [722] & !i[1817]) | ( l_40 [723] &  i[1817]);
assign l_39[371]    = ( l_40 [724] & !i[1817]) | ( l_40 [725] &  i[1817]);
assign l_39[372]    = ( l_40 [726] & !i[1817]) | ( l_40 [727] &  i[1817]);
assign l_39[373]    = ( l_40 [728] & !i[1817]) | ( l_40 [729] &  i[1817]);
assign l_39[374]    = ( l_40 [730] & !i[1817]) | ( l_40 [731] &  i[1817]);
assign l_39[375]    = ( l_40 [732] & !i[1817]) | ( l_40 [733] &  i[1817]);
assign l_39[376]    = ( l_40 [734] & !i[1817]) | ( l_40 [735] &  i[1817]);
assign l_39[377]    = ( l_40 [736] & !i[1817]) | ( l_40 [737] &  i[1817]);
assign l_39[378]    = ( l_40 [738] & !i[1817]) | ( l_40 [739] &  i[1817]);
assign l_39[379]    = ( l_40 [740] & !i[1817]) | ( l_40 [741] &  i[1817]);
assign l_39[380]    = ( l_40 [742] & !i[1817]) | ( l_40 [743] &  i[1817]);
assign l_39[381]    = ( l_40 [744] & !i[1817]) | ( l_40 [745] &  i[1817]);
assign l_39[382]    = ( l_40 [746] & !i[1817]) | ( l_40 [747] &  i[1817]);
assign l_39[383]    = ( l_40 [748] & !i[1817]) | ( l_40 [749] &  i[1817]);
assign l_39[384]    = ( l_40 [750] & !i[1817]) | ( l_40 [751] &  i[1817]);
assign l_39[385]    = ( l_40 [752] & !i[1817]) | ( l_40 [753] &  i[1817]);
assign l_39[386]    = ( l_40 [754] & !i[1817]) | ( l_40 [755] &  i[1817]);
assign l_39[387]    = ( l_40 [756] & !i[1817]) | ( l_40 [757] &  i[1817]);
assign l_39[388]    = ( l_40 [758] & !i[1817]) | ( l_40 [759] &  i[1817]);
assign l_39[389]    = ( l_40 [760] & !i[1817]) | ( l_40 [761] &  i[1817]);
assign l_39[390]    = ( l_40 [762] & !i[1817]) | ( l_40 [763] &  i[1817]);
assign l_39[391]    = ( l_40 [764] & !i[1817]) | ( l_40 [765] &  i[1817]);
assign l_39[392]    = ( l_40 [766] & !i[1817]) | ( l_40 [767] &  i[1817]);
assign l_39[393]    = ( l_40 [768] & !i[1817]) | ( l_40 [769] &  i[1817]);
assign l_39[394]    = ( l_40 [770] & !i[1817]) | ( l_40 [771] &  i[1817]);
assign l_39[395]    = ( l_40 [772] & !i[1817]) | ( l_40 [773] &  i[1817]);
assign l_39[396]    = ( l_40 [774] & !i[1817]) | ( l_40 [775] &  i[1817]);
assign l_39[397]    = ( l_40 [776] & !i[1817]) | ( l_40 [777] &  i[1817]);
assign l_39[398]    = ( l_40 [778] & !i[1817]) | ( l_40 [779] &  i[1817]);
assign l_39[399]    = ( l_40 [780] & !i[1817]) | ( l_40 [781] &  i[1817]);
assign l_39[400]    = ( l_40 [782] & !i[1817]) | ( l_40 [783] &  i[1817]);
assign l_39[401]    = ( l_40 [784] & !i[1817]) | ( l_40 [785] &  i[1817]);
assign l_39[402]    = ( l_40 [786] & !i[1817]) | ( l_40 [787] &  i[1817]);
assign l_39[403]    = ( l_40 [788] & !i[1817]) | ( l_40 [789] &  i[1817]);
assign l_39[404]    = ( l_40 [790] & !i[1817]) | ( l_40 [791] &  i[1817]);
assign l_39[405]    = ( l_40 [792] & !i[1817]) | ( l_40 [793] &  i[1817]);
assign l_39[406]    = ( l_40 [794] & !i[1817]) | ( l_40 [795] &  i[1817]);
assign l_39[407]    = ( l_40 [796] & !i[1817]) | ( l_40 [797] &  i[1817]);
assign l_39[408]    = ( l_40 [798] & !i[1817]) | ( l_40 [799] &  i[1817]);
assign l_39[409]    = ( l_40 [800] & !i[1817]) | ( l_40 [801] &  i[1817]);
assign l_39[410]    = ( l_40 [802] & !i[1817]) | ( l_40 [803] &  i[1817]);
assign l_39[411]    = ( l_40 [804] & !i[1817]) | ( l_40 [805] &  i[1817]);
assign l_39[412]    = ( l_40 [806] & !i[1817]) | ( l_40 [807] &  i[1817]);
assign l_39[413]    = ( l_40 [808] & !i[1817]) | ( l_40 [809] &  i[1817]);
assign l_39[414]    = ( l_40 [810] & !i[1817]) | ( l_40 [811] &  i[1817]);
assign l_39[415]    = ( l_40 [812] & !i[1817]) | ( l_40 [813] &  i[1817]);
assign l_39[416]    = ( l_40 [814] & !i[1817]) | ( l_40 [815] &  i[1817]);
assign l_39[417]    = ( l_40 [816] & !i[1817]) | ( l_40 [817] &  i[1817]);
assign l_39[418]    = ( l_40 [818] & !i[1817]) | ( l_40 [819] &  i[1817]);
assign l_39[419]    = ( l_40 [820] & !i[1817]) | ( l_40 [821] &  i[1817]);
assign l_39[420]    = ( l_40 [822] & !i[1817]) | ( l_40 [823] &  i[1817]);
assign l_39[421]    = ( l_40 [824] & !i[1817]) | ( l_40 [825] &  i[1817]);
assign l_39[422]    = ( l_40 [826] & !i[1817]) | ( l_40 [827] &  i[1817]);
assign l_39[423]    = ( l_40 [828] & !i[1817]) | ( l_40 [829] &  i[1817]);
assign l_39[424]    = ( l_40 [830] & !i[1817]) | ( l_40 [831] &  i[1817]);
assign l_39[425]    = ( l_40 [832] & !i[1817]) | ( l_40 [833] &  i[1817]);
assign l_39[426]    = ( l_40 [834] & !i[1817]) | ( l_40 [835] &  i[1817]);
assign l_39[427]    = ( l_40 [836] & !i[1817]) | ( l_40 [837] &  i[1817]);
assign l_39[428]    = ( l_40 [838] & !i[1817]) | ( l_40 [839] &  i[1817]);
assign l_39[429]    = ( l_40 [840] & !i[1817]) | ( l_40 [841] &  i[1817]);
assign l_39[430]    = ( l_40 [842] & !i[1817]) | ( l_40 [843] &  i[1817]);
assign l_39[431]    = ( l_40 [844] & !i[1817]) | ( l_40 [845] &  i[1817]);
assign l_39[432]    = ( l_40 [846] & !i[1817]) | ( l_40 [847] &  i[1817]);
assign l_39[433]    = ( l_40 [848] & !i[1817]) | ( l_40 [849] &  i[1817]);
assign l_39[434]    = ( l_40 [850] & !i[1817]) | ( l_40 [851] &  i[1817]);
assign l_39[435]    = ( l_40 [852] & !i[1817]) | ( l_40 [853] &  i[1817]);
assign l_39[436]    = ( l_40 [854] & !i[1817]) | ( l_40 [855] &  i[1817]);
assign l_39[437]    = ( l_40 [856] & !i[1817]) | ( l_40 [857] &  i[1817]);
assign l_39[438]    = ( l_40 [858] & !i[1817]) | ( l_40 [859] &  i[1817]);
assign l_39[439]    = ( l_40 [860] & !i[1817]) | ( l_40 [861] &  i[1817]);
assign l_39[440]    = ( l_40 [862] & !i[1817]) | ( l_40 [863] &  i[1817]);
assign l_39[441]    = ( l_40 [864] & !i[1817]) | ( l_40 [865] &  i[1817]);
assign l_39[442]    = ( l_40 [866] & !i[1817]) | ( l_40 [867] &  i[1817]);
assign l_39[443]    = ( l_40 [868] & !i[1817]) | ( l_40 [869] &  i[1817]);
assign l_39[444]    = ( l_40 [870] & !i[1817]) | ( l_40 [871] &  i[1817]);
assign l_39[445]    = ( l_40 [872] & !i[1817]) | ( l_40 [873] &  i[1817]);
assign l_39[446]    = ( l_40 [874] & !i[1817]) | ( l_40 [875] &  i[1817]);
assign l_39[447]    = ( l_40 [876] & !i[1817]) | ( l_40 [877] &  i[1817]);
assign l_39[448]    = ( l_40 [878] & !i[1817]) | ( l_40 [879] &  i[1817]);
assign l_39[449]    = ( l_40 [880] & !i[1817]) | ( l_40 [881] &  i[1817]);
assign l_39[450]    = ( l_40 [882] & !i[1817]) | ( l_40 [883] &  i[1817]);
assign l_39[451]    = ( l_40 [884] & !i[1817]) | ( l_40 [885] &  i[1817]);
assign l_39[452]    = ( l_40 [886] & !i[1817]) | ( l_40 [887] &  i[1817]);
assign l_39[453]    = ( l_40 [888] & !i[1817]) | ( l_40 [889] &  i[1817]);
assign l_39[454]    = ( l_40 [890] & !i[1817]) | ( l_40 [891] &  i[1817]);
assign l_39[455]    = ( l_40 [892] & !i[1817]) | ( l_40 [893] &  i[1817]);
assign l_39[456]    = ( l_40 [894] & !i[1817]) | ( l_40 [895] &  i[1817]);
assign l_39[457]    = ( l_40 [896] & !i[1817]) | ( l_40 [897] &  i[1817]);
assign l_39[458]    = ( l_40 [898] & !i[1817]) | ( l_40 [899] &  i[1817]);
assign l_39[459]    = ( l_40 [900] & !i[1817]) | ( l_40 [901] &  i[1817]);
assign l_39[460]    = ( l_40 [902] & !i[1817]) | ( l_40 [903] &  i[1817]);
assign l_39[461]    = ( l_40 [904] & !i[1817]) | ( l_40 [905] &  i[1817]);
assign l_39[462]    = ( l_40 [906] & !i[1817]) | ( l_40 [907] &  i[1817]);
assign l_39[463]    = ( l_40 [908] & !i[1817]) | ( l_40 [909] &  i[1817]);
assign l_39[464]    = ( l_40 [910] & !i[1817]) | ( l_40 [911] &  i[1817]);
assign l_39[465]    = ( l_40 [912] & !i[1817]) | ( l_40 [913] &  i[1817]);
assign l_39[466]    = ( l_40 [914] & !i[1817]) | ( l_40 [915] &  i[1817]);
assign l_39[467]    = ( l_40 [916] & !i[1817]) | ( l_40 [917] &  i[1817]);
assign l_39[468]    = ( l_40 [918] & !i[1817]) | ( l_40 [919] &  i[1817]);
assign l_39[469]    = ( l_40 [920] & !i[1817]) | ( l_40 [921] &  i[1817]);
assign l_39[470]    = ( l_40 [922] & !i[1817]) | ( l_40 [923] &  i[1817]);
assign l_39[471]    = ( l_40 [924] & !i[1817]) | ( l_40 [925] &  i[1817]);
assign l_39[472]    = ( l_40 [926] & !i[1817]) | ( l_40 [927] &  i[1817]);
assign l_39[473]    = ( l_40 [928] & !i[1817]) | ( l_40 [929] &  i[1817]);
assign l_39[474]    = ( l_40 [930] & !i[1817]) | ( l_40 [931] &  i[1817]);
assign l_39[475]    = ( l_40 [932] & !i[1817]) | ( l_40 [933] &  i[1817]);
assign l_39[476]    = ( l_40 [934] & !i[1817]) | ( l_40 [935] &  i[1817]);
assign l_39[477]    = ( l_40 [936] & !i[1817]) | ( l_40 [937] &  i[1817]);
assign l_39[478]    = ( l_40 [938] & !i[1817]) | ( l_40 [939] &  i[1817]);
assign l_39[479]    = ( l_40 [940] & !i[1817]) | ( l_40 [941] &  i[1817]);
assign l_39[480]    = ( l_40 [942] & !i[1817]) | ( l_40 [943] &  i[1817]);
assign l_39[481]    = ( l_40 [944] & !i[1817]) | ( l_40 [945] &  i[1817]);
assign l_39[482]    = ( l_40 [946] & !i[1817]) | ( l_40 [947] &  i[1817]);
assign l_39[483]    = ( l_40 [948] & !i[1817]) | ( l_40 [949] &  i[1817]);
assign l_39[484]    = ( l_40 [950] & !i[1817]) | ( l_40 [951] &  i[1817]);
assign l_39[485]    = ( l_40 [952] & !i[1817]) | ( l_40 [953] &  i[1817]);
assign l_39[486]    = ( l_40 [954] & !i[1817]) | ( l_40 [955] &  i[1817]);
assign l_39[487]    = ( l_40 [956] & !i[1817]) | ( l_40 [957] &  i[1817]);
assign l_39[488]    = ( l_40 [958] & !i[1817]) | ( l_40 [959] &  i[1817]);
assign l_39[489]    = ( l_40 [960] & !i[1817]) | ( l_40 [961] &  i[1817]);
assign l_39[490]    = ( l_40 [962] & !i[1817]) | ( l_40 [963] &  i[1817]);
assign l_39[491]    = ( l_40 [964] & !i[1817]) | ( l_40 [965] &  i[1817]);
assign l_39[492]    = ( l_40 [966] & !i[1817]) | ( l_40 [967] &  i[1817]);
assign l_39[493]    = ( l_40 [968] & !i[1817]) | ( l_40 [969] &  i[1817]);
assign l_39[494]    = ( l_40 [970] & !i[1817]) | ( l_40 [971] &  i[1817]);
assign l_39[495]    = ( l_40 [972] & !i[1817]) | ( l_40 [973] &  i[1817]);
assign l_39[496]    = ( l_40 [974] & !i[1817]) | ( l_40 [975] &  i[1817]);
assign l_39[497]    = ( l_40 [976] & !i[1817]) | ( l_40 [977] &  i[1817]);
assign l_39[498]    = ( l_40 [978] & !i[1817]) | ( l_40 [979] &  i[1817]);
assign l_39[499]    = ( l_40 [980] & !i[1817]) | ( l_40 [981] &  i[1817]);
assign l_39[500]    = ( l_40 [982] & !i[1817]) | ( l_40 [983] &  i[1817]);
assign l_39[501]    = ( l_40 [984] & !i[1817]) | ( l_40 [985] &  i[1817]);
assign l_39[502]    = ( l_40 [986] & !i[1817]) | ( l_40 [987] &  i[1817]);
assign l_39[503]    = ( l_40 [988] & !i[1817]) | ( l_40 [989] &  i[1817]);
assign l_39[504]    = ( l_40 [990] & !i[1817]) | ( l_40 [991] &  i[1817]);
assign l_39[505]    = ( l_40 [992] & !i[1817]) | ( l_40 [993] &  i[1817]);
assign l_39[506]    = ( l_40 [994] & !i[1817]) | ( l_40 [995] &  i[1817]);
assign l_39[507]    = ( l_40 [996] & !i[1817]) | ( l_40 [997] &  i[1817]);
assign l_39[508]    = ( l_40 [998] & !i[1817]) | ( l_40 [999] &  i[1817]);
assign l_39[509]    = ( l_40 [1000] & !i[1817]) | ( l_40 [1001] &  i[1817]);
assign l_39[510]    = ( l_40 [1002] & !i[1817]) | ( l_40 [1003] &  i[1817]);
assign l_39[511]    = ( l_40 [1004] & !i[1817]) | ( l_40 [1005] &  i[1817]);
assign l_39[512]    = ( l_40 [1006] & !i[1817]) | ( l_40 [1007] &  i[1817]);
assign l_39[513]    = ( l_40 [1008] & !i[1817]) | ( l_40 [1009] &  i[1817]);
assign l_39[514]    = ( l_40 [1010] & !i[1817]) | ( l_40 [1011] &  i[1817]);
assign l_39[515]    = ( l_40 [1012] & !i[1817]) | ( l_40 [1013] &  i[1817]);
assign l_39[516]    = ( l_40 [1014] & !i[1817]) | ( l_40 [1015] &  i[1817]);
assign l_39[517]    = ( l_40 [1016] & !i[1817]) | ( l_40 [1017] &  i[1817]);
assign l_39[518]    = ( l_40 [1018] & !i[1817]) | ( l_40 [1019] &  i[1817]);
assign l_39[519]    = ( l_40 [1020] & !i[1817]) | ( l_40 [1021] &  i[1817]);
assign l_39[520]    = ( l_40 [1022] & !i[1817]) | ( l_40 [1023] &  i[1817]);
assign l_39[521]    = ( l_40 [1024] & !i[1817]) | ( l_40 [1025] &  i[1817]);
assign l_39[522]    = ( l_40 [1026] & !i[1817]) | ( l_40 [1027] &  i[1817]);
assign l_39[523]    = ( l_40 [1028] & !i[1817]) | ( l_40 [1029] &  i[1817]);
assign l_39[524]    = ( l_40 [1030] & !i[1817]) | ( l_40 [1031] &  i[1817]);
assign l_39[525]    = ( l_40 [1032] & !i[1817]) | ( l_40 [1033] &  i[1817]);
assign l_39[526]    = ( l_40 [1034] & !i[1817]) | ( l_40 [1035] &  i[1817]);
assign l_39[527]    = ( l_40 [1036] & !i[1817]) | ( l_40 [1037] &  i[1817]);
assign l_39[528]    = ( l_40 [1038] & !i[1817]) | ( l_40 [1039] &  i[1817]);
assign l_39[529]    = ( l_40 [1040] & !i[1817]) | ( l_40 [1041] &  i[1817]);
assign l_39[530]    = ( l_40 [1042] & !i[1817]) | ( l_40 [1043] &  i[1817]);
assign l_39[531]    = ( l_40 [1044] & !i[1817]) | ( l_40 [1045] &  i[1817]);
assign l_39[532]    = ( l_40 [1046] & !i[1817]) | ( l_40 [1047] &  i[1817]);
assign l_39[533]    = ( l_40 [1048] & !i[1817]) | ( l_40 [1049] &  i[1817]);
assign l_39[534]    = ( l_40 [1050] & !i[1817]) | ( l_40 [1051] &  i[1817]);
assign l_39[535]    = ( l_40 [1052] & !i[1817]) | ( l_40 [1053] &  i[1817]);
assign l_39[536]    = ( l_40 [1054] & !i[1817]) | ( l_40 [1055] &  i[1817]);
assign l_39[537]    = ( l_40 [1056] & !i[1817]) | ( l_40 [1057] &  i[1817]);
assign l_39[538]    = ( l_40 [1058] & !i[1817]) | ( l_40 [1059] &  i[1817]);
assign l_39[539]    = ( l_40 [1060] & !i[1817]) | ( l_40 [1061] &  i[1817]);
assign l_39[540]    = ( l_40 [1062] & !i[1817]) | ( l_40 [1063] &  i[1817]);
assign l_39[541]    = ( l_40 [1064] & !i[1817]) | ( l_40 [1065] &  i[1817]);
assign l_39[542]    = ( l_40 [1066] & !i[1817]) | ( l_40 [1067] &  i[1817]);
assign l_39[543]    = ( l_40 [1068] & !i[1817]) | ( l_40 [1069] &  i[1817]);
assign l_39[544]    = ( l_40 [1070] & !i[1817]) | ( l_40 [1071] &  i[1817]);
assign l_39[545]    = ( l_40 [1072] & !i[1817]) | ( l_40 [1073] &  i[1817]);
assign l_39[546]    = ( l_40 [1074] & !i[1817]) | ( l_40 [1075] &  i[1817]);
assign l_39[547]    = ( l_40 [1076] & !i[1817]) | ( l_40 [1077] &  i[1817]);
assign l_39[548]    = ( l_40 [1078] & !i[1817]) | ( l_40 [1079] &  i[1817]);
assign l_39[549]    = ( l_40 [1080] & !i[1817]) | ( l_40 [1081] &  i[1817]);
assign l_39[550]    = ( l_40 [1082] & !i[1817]) | ( l_40 [1083] &  i[1817]);
assign l_39[551]    = ( l_40 [1084] & !i[1817]) | ( l_40 [1085] &  i[1817]);
assign l_39[552]    = ( l_40 [1086] & !i[1817]) | ( l_40 [1087] &  i[1817]);
assign l_39[553]    = ( l_40 [1088] & !i[1817]) | ( l_40 [1089] &  i[1817]);
assign l_39[554]    = ( l_40 [1090] & !i[1817]) | ( l_40 [1091] &  i[1817]);
assign l_39[555]    = ( l_40 [1092] & !i[1817]) | ( l_40 [1093] &  i[1817]);
assign l_39[556]    = ( l_40 [1094] & !i[1817]) | ( l_40 [1095] &  i[1817]);
assign l_39[557]    = ( l_40 [1096] & !i[1817]) | ( l_40 [1097] &  i[1817]);
assign l_39[558]    = ( l_40 [1098] & !i[1817]) | ( l_40 [1099] &  i[1817]);
assign l_39[559]    = ( l_40 [1100] & !i[1817]) | ( l_40 [1101] &  i[1817]);
assign l_39[560]    = ( l_40 [1102] & !i[1817]) | ( l_40 [1103] &  i[1817]);
assign l_39[561]    = ( l_40 [1104] & !i[1817]) | ( l_40 [1105] &  i[1817]);
assign l_39[562]    = ( l_40 [1106] & !i[1817]) | ( l_40 [1107] &  i[1817]);
assign l_39[563]    = ( l_40 [1108] & !i[1817]) | ( l_40 [1109] &  i[1817]);
assign l_39[564]    = ( l_40 [1110] & !i[1817]) | ( l_40 [1111] &  i[1817]);
assign l_39[565]    = ( l_40 [1112] & !i[1817]) | ( l_40 [1113] &  i[1817]);
assign l_39[566]    = ( l_40 [1114] & !i[1817]) | ( l_40 [1115] &  i[1817]);
assign l_39[567]    = ( l_40 [1116] & !i[1817]) | ( l_40 [1117] &  i[1817]);
assign l_39[568]    = ( l_40 [1118] & !i[1817]) | ( l_40 [1119] &  i[1817]);
assign l_39[569]    = ( l_40 [1120] & !i[1817]) | ( l_40 [1121] &  i[1817]);
assign l_39[570]    = ( l_40 [1122] & !i[1817]) | ( l_40 [1123] &  i[1817]);
assign l_39[571]    = ( l_40 [1124] & !i[1817]) | ( l_40 [1125] &  i[1817]);
assign l_39[572]    = ( l_40 [1126] & !i[1817]) | ( l_40 [1127] &  i[1817]);
assign l_39[573]    = ( l_40 [1128] & !i[1817]) | ( l_40 [1129] &  i[1817]);
assign l_39[574]    = ( l_40 [1130] & !i[1817]) | ( l_40 [1131] &  i[1817]);
assign l_39[575]    = ( l_40 [1132] & !i[1817]) | ( l_40 [1133] &  i[1817]);
assign l_39[576]    = ( l_40 [1134] & !i[1817]) | ( l_40 [1135] &  i[1817]);
assign l_39[577]    = ( l_40 [1136] & !i[1817]) | ( l_40 [1137] &  i[1817]);
assign l_39[578]    = ( l_40 [1138] & !i[1817]) | ( l_40 [1139] &  i[1817]);
assign l_39[579]    = ( l_40 [1140] & !i[1817]) | ( l_40 [1141] &  i[1817]);
assign l_39[580]    = ( l_40 [1142] & !i[1817]) | ( l_40 [1143] &  i[1817]);
assign l_39[581]    = ( l_40 [1144] & !i[1817]) | ( l_40 [1145] &  i[1817]);
assign l_39[582]    = ( l_40 [1146] & !i[1817]) | ( l_40 [1147] &  i[1817]);
assign l_39[583]    = ( l_40 [1148] & !i[1817]) | ( l_40 [1149] &  i[1817]);
assign l_39[584]    = ( l_40 [1150] & !i[1817]) | ( l_40 [1151] &  i[1817]);
assign l_39[585]    = ( l_40 [1152] & !i[1817]) | ( l_40 [1153] &  i[1817]);
assign l_39[586]    = ( l_40 [1154] & !i[1817]) | ( l_40 [1155] &  i[1817]);
assign l_39[587]    = ( l_40 [1156] & !i[1817]) | ( l_40 [1157] &  i[1817]);
assign l_39[588]    = ( l_40 [1158] & !i[1817]) | ( l_40 [1159] &  i[1817]);
assign l_39[589]    = ( l_40 [1160] & !i[1817]) | ( l_40 [1161] &  i[1817]);
assign l_39[590]    = ( l_40 [1162] & !i[1817]) | ( l_40 [1163] &  i[1817]);
assign l_39[591]    = ( l_40 [1164] & !i[1817]) | ( l_40 [1165] &  i[1817]);
assign l_39[592]    = ( l_40 [1166] & !i[1817]) | ( l_40 [1167] &  i[1817]);
assign l_39[593]    = ( l_40 [1168] & !i[1817]) | ( l_40 [1169] &  i[1817]);
assign l_39[594]    = ( l_40 [1170] & !i[1817]) | ( l_40 [1171] &  i[1817]);
assign l_39[595]    = ( l_40 [1172] & !i[1817]) | ( l_40 [1173] &  i[1817]);
assign l_39[596]    = ( l_40 [1174] & !i[1817]) | ( l_40 [1175] &  i[1817]);
assign l_39[597]    = ( l_40 [1176] & !i[1817]) | ( l_40 [1177] &  i[1817]);
assign l_39[598]    = ( l_40 [1178] & !i[1817]) | ( l_40 [1179] &  i[1817]);
assign l_39[599]    = ( l_40 [1180] & !i[1817]) | ( l_40 [1181] &  i[1817]);
assign l_39[600]    = ( l_40 [1182] & !i[1817]) | ( l_40 [1183] &  i[1817]);
assign l_39[601]    = ( l_40 [1184] & !i[1817]) | ( l_40 [1185] &  i[1817]);
assign l_39[602]    = ( l_40 [1186] & !i[1817]) | ( l_40 [1187] &  i[1817]);
assign l_39[603]    = ( l_40 [1188] & !i[1817]) | ( l_40 [1189] &  i[1817]);
assign l_39[604]    = ( l_40 [1190] & !i[1817]) | ( l_40 [1191] &  i[1817]);
assign l_39[605]    = ( l_40 [1192] & !i[1817]) | ( l_40 [1193] &  i[1817]);
assign l_39[606]    = ( l_40 [1194] & !i[1817]) | ( l_40 [1195] &  i[1817]);
assign l_39[607]    = ( l_40 [1196] & !i[1817]) | ( l_40 [1197] &  i[1817]);
assign l_39[608]    = ( l_40 [1198] & !i[1817]) | ( l_40 [1199] &  i[1817]);
assign l_39[609]    = ( l_40 [1200] & !i[1817]) | ( l_40 [1201] &  i[1817]);
assign l_39[610]    = ( l_40 [1202] & !i[1817]) | ( l_40 [1203] &  i[1817]);
assign l_39[611]    = ( l_40 [1204] & !i[1817]) | ( l_40 [1205] &  i[1817]);
assign l_39[612]    = ( l_40 [1206] & !i[1817]) | ( l_40 [1207] &  i[1817]);
assign l_39[613]    = ( l_40 [1208] & !i[1817]) | ( l_40 [1209] &  i[1817]);
assign l_39[614]    = ( l_40 [1210] & !i[1817]) | ( l_40 [1211] &  i[1817]);
assign l_39[615]    = ( l_40 [1212] & !i[1817]) | ( l_40 [1213] &  i[1817]);
assign l_39[616]    = ( l_40 [1214] & !i[1817]) | ( l_40 [1215] &  i[1817]);
assign l_39[617]    = ( l_40 [1216] & !i[1817]) | ( l_40 [1217] &  i[1817]);
assign l_39[618]    = ( l_40 [1218] & !i[1817]) | ( l_40 [1219] &  i[1817]);
assign l_39[619]    = ( l_40 [1220] & !i[1817]) | ( l_40 [1221] &  i[1817]);
assign l_39[620]    = ( l_40 [1222] & !i[1817]) | ( l_40 [1223] &  i[1817]);
assign l_39[621]    = ( l_40 [1224] & !i[1817]) | ( l_40 [1225] &  i[1817]);
assign l_39[622]    = ( l_40 [1226] & !i[1817]) | ( l_40 [1227] &  i[1817]);
assign l_39[623]    = ( l_40 [1228] & !i[1817]) | ( l_40 [1229] &  i[1817]);
assign l_39[624]    = ( l_40 [1230] & !i[1817]) | ( l_40 [1231] &  i[1817]);
assign l_39[625]    = ( l_40 [1232] & !i[1817]) | ( l_40 [1233] &  i[1817]);
assign l_39[626]    = ( l_40 [1234] & !i[1817]) | ( l_40 [1235] &  i[1817]);
assign l_39[627]    = ( l_40 [1236] & !i[1817]) | ( l_40 [1237] &  i[1817]);
assign l_39[628]    = ( l_40 [1238] & !i[1817]) | ( l_40 [1239] &  i[1817]);
assign l_39[629]    = ( l_40 [1240] & !i[1817]) | ( l_40 [1241] &  i[1817]);
assign l_39[630]    = ( l_40 [1242] & !i[1817]) | ( l_40 [1243] &  i[1817]);
assign l_39[631]    = ( l_40 [1244] & !i[1817]) | ( l_40 [1245] &  i[1817]);
assign l_39[632]    = ( l_40 [1246] & !i[1817]) | ( l_40 [1247] &  i[1817]);
assign l_39[633]    = ( l_40 [1248] & !i[1817]) | ( l_40 [1249] &  i[1817]);
assign l_39[634]    = ( l_40 [1250] & !i[1817]) | ( l_40 [1251] &  i[1817]);
assign l_39[635]    = ( l_40 [1252] & !i[1817]) | ( l_40 [1253] &  i[1817]);
assign l_39[636]    = ( l_40 [1254] & !i[1817]) | ( l_40 [1255] &  i[1817]);
assign l_39[637]    = ( l_40 [1256] & !i[1817]) | ( l_40 [1257] &  i[1817]);
assign l_39[638]    = ( l_40 [1258] & !i[1817]) | ( l_40 [1259] &  i[1817]);
assign l_39[639]    = ( l_40 [1260] & !i[1817]) | ( l_40 [1261] &  i[1817]);
assign l_39[640]    = ( l_40 [1262] & !i[1817]) | ( l_40 [1263] &  i[1817]);
assign l_39[641]    = ( l_40 [1264] & !i[1817]) | ( l_40 [1265] &  i[1817]);
assign l_39[642]    = ( l_40 [1266] & !i[1817]) | ( l_40 [1267] &  i[1817]);
assign l_39[643]    = ( l_40 [1268] & !i[1817]) | ( l_40 [1269] &  i[1817]);
assign l_39[644]    = ( l_40 [1270] & !i[1817]) | ( l_40 [1271] &  i[1817]);
assign l_39[645]    = ( l_40 [1272] & !i[1817]) | ( l_40 [1273] &  i[1817]);
assign l_39[646]    = ( l_40 [1274] & !i[1817]) | ( l_40 [1275] &  i[1817]);
assign l_39[647]    = ( l_40 [1276] & !i[1817]) | ( l_40 [1277] &  i[1817]);
assign l_39[648]    = ( l_40 [1278] & !i[1817]) | ( l_40 [1279] &  i[1817]);
assign l_39[649]    = ( l_40 [1280] & !i[1817]) | ( l_40 [1281] &  i[1817]);
assign l_39[650]    = ( l_40 [1282] & !i[1817]) | ( l_40 [1283] &  i[1817]);
assign l_39[651]    = ( l_40 [1284] & !i[1817]) | ( l_40 [1285] &  i[1817]);
assign l_39[652]    = ( l_40 [1286] & !i[1817]) | ( l_40 [1287] &  i[1817]);
assign l_39[653]    = ( l_40 [1288] & !i[1817]) | ( l_40 [1289] &  i[1817]);
assign l_39[654]    = ( l_40 [1290] & !i[1817]) | ( l_40 [1291] &  i[1817]);
assign l_39[655]    = ( l_40 [1292] & !i[1817]) | ( l_40 [1293] &  i[1817]);
assign l_39[656]    = ( l_40 [1294] & !i[1817]) | ( l_40 [1295] &  i[1817]);
assign l_39[657]    = ( l_40 [1296] & !i[1817]) | ( l_40 [1297] &  i[1817]);
assign l_39[658]    = ( l_40 [1298] & !i[1817]) | ( l_40 [1299] &  i[1817]);
assign l_39[659]    = ( l_40 [1300] & !i[1817]) | ( l_40 [1301] &  i[1817]);
assign l_39[660]    = ( l_40 [1302] & !i[1817]) | ( l_40 [1303] &  i[1817]);
assign l_39[661]    = ( l_40 [1304] & !i[1817]) | ( l_40 [1305] &  i[1817]);
assign l_39[662]    = ( l_40 [1306] & !i[1817]) | ( l_40 [1307] &  i[1817]);
assign l_39[663]    = ( l_40 [1308] & !i[1817]) | ( l_40 [1309] &  i[1817]);
assign l_39[664]    = ( l_40 [1310] & !i[1817]) | ( l_40 [1311] &  i[1817]);
assign l_39[665]    = ( l_40 [1312] & !i[1817]) | ( l_40 [1313] &  i[1817]);
assign l_39[666]    = ( l_40 [1314] & !i[1817]) | ( l_40 [1315] &  i[1817]);
assign l_39[667]    = ( l_40 [1316] & !i[1817]) | ( l_40 [1317] &  i[1817]);
assign l_39[668]    = ( l_40 [1318] & !i[1817]) | ( l_40 [1319] &  i[1817]);
assign l_39[669]    = ( l_40 [1320] & !i[1817]) | ( l_40 [1321] &  i[1817]);
assign l_39[670]    = ( l_40 [1322] & !i[1817]) | ( l_40 [1323] &  i[1817]);
assign l_39[671]    = ( l_40 [1324] & !i[1817]) | ( l_40 [1325] &  i[1817]);
assign l_39[672]    = ( l_40 [1326] & !i[1817]) | ( l_40 [1327] &  i[1817]);
assign l_39[673]    = ( l_40 [1328] & !i[1817]) | ( l_40 [1329] &  i[1817]);
assign l_39[674]    = ( l_40 [1330] & !i[1817]) | ( l_40 [1331] &  i[1817]);
assign l_39[675]    = ( l_40 [1332] & !i[1817]) | ( l_40 [1333] &  i[1817]);
assign l_39[676]    = ( l_40 [1334] & !i[1817]) | ( l_40 [1335] &  i[1817]);
assign l_39[677]    = ( l_40 [1336] & !i[1817]) | ( l_40 [1337] &  i[1817]);
assign l_39[678]    = ( l_40 [1338] & !i[1817]) | ( l_40 [1339] &  i[1817]);
assign l_39[679]    = ( l_40 [1340] & !i[1817]) | ( l_40 [1341] &  i[1817]);
assign l_39[680]    = ( l_40 [1342] & !i[1817]) | ( l_40 [1343] &  i[1817]);
assign l_39[681]    = ( l_40 [1344] & !i[1817]) | ( l_40 [1345] &  i[1817]);
assign l_39[682]    = ( l_40 [1346] & !i[1817]) | ( l_40 [1347] &  i[1817]);
assign l_39[683]    = ( l_40 [1348] & !i[1817]) | ( l_40 [1349] &  i[1817]);
assign l_39[684]    = ( l_40 [1350] & !i[1817]) | ( l_40 [1351] &  i[1817]);
assign l_39[685]    = ( l_40 [1352] & !i[1817]) | ( l_40 [1353] &  i[1817]);
assign l_39[686]    = ( l_40 [1354] & !i[1817]) | ( l_40 [1355] &  i[1817]);
assign l_39[687]    = ( l_40 [1356] & !i[1817]) | ( l_40 [1357] &  i[1817]);
assign l_39[688]    = ( l_40 [1358] & !i[1817]) | ( l_40 [1359] &  i[1817]);
assign l_39[689]    = ( l_40 [1360] & !i[1817]) | ( l_40 [1361] &  i[1817]);
assign l_39[690]    = ( l_40 [1362] & !i[1817]) | ( l_40 [1363] &  i[1817]);
assign l_39[691]    = ( l_40 [1364] & !i[1817]) | ( l_40 [1365] &  i[1817]);
assign l_39[692]    = ( l_40 [1366] & !i[1817]) | ( l_40 [1367] &  i[1817]);
assign l_39[693]    = ( l_40 [1368] & !i[1817]) | ( l_40 [1369] &  i[1817]);
assign l_39[694]    = ( l_40 [1370] & !i[1817]) | ( l_40 [1371] &  i[1817]);
assign l_39[695]    = ( l_40 [1372] & !i[1817]) | ( l_40 [1373] &  i[1817]);
assign l_39[696]    = ( l_40 [1374] & !i[1817]) | ( l_40 [1375] &  i[1817]);
assign l_39[697]    = ( l_40 [1376] & !i[1817]) | ( l_40 [1377] &  i[1817]);
assign l_39[698]    = ( l_40 [1378] & !i[1817]) | ( l_40 [1379] &  i[1817]);
assign l_39[699]    = ( l_40 [1380] & !i[1817]) | ( l_40 [1381] &  i[1817]);
assign l_39[700]    = ( l_40 [1382] & !i[1817]) | ( l_40 [1383] &  i[1817]);
assign l_39[701]    = ( l_40 [1384] & !i[1817]) | ( l_40 [1385] &  i[1817]);
assign l_39[702]    = ( l_40 [1386] & !i[1817]) | ( l_40 [1387] &  i[1817]);
assign l_39[703]    = ( l_40 [1388] & !i[1817]) | ( l_40 [1389] &  i[1817]);
assign l_39[704]    = ( l_40 [1390] & !i[1817]) | ( l_40 [1391] &  i[1817]);
assign l_39[705]    = ( l_40 [1392] & !i[1817]) | ( l_40 [1393] &  i[1817]);
assign l_39[706]    = ( l_40 [1394] & !i[1817]) | ( l_40 [1395] &  i[1817]);
assign l_39[707]    = ( l_40 [1396] & !i[1817]) | ( l_40 [1397] &  i[1817]);
assign l_39[708]    = ( l_40 [1398] & !i[1817]) | ( l_40 [1399] &  i[1817]);
assign l_39[709]    = ( l_40 [1400] & !i[1817]) | ( l_40 [1401] &  i[1817]);
assign l_39[710]    = ( l_40 [1402] & !i[1817]) | ( l_40 [1403] &  i[1817]);
assign l_39[711]    = ( l_40 [1404] & !i[1817]) | ( l_40 [1405] &  i[1817]);
assign l_39[712]    = ( l_40 [1406] & !i[1817]) | ( l_40 [1407] &  i[1817]);
assign l_39[713]    = ( l_40 [1408] & !i[1817]) | ( l_40 [1409] &  i[1817]);
assign l_39[714]    = ( l_40 [1410] & !i[1817]) | ( l_40 [1411] &  i[1817]);
assign l_39[715]    = ( l_40 [1412] & !i[1817]) | ( l_40 [1413] &  i[1817]);
assign l_39[716]    = ( l_40 [1414] & !i[1817]) | ( l_40 [1415] &  i[1817]);
assign l_39[717]    = ( l_40 [1416] & !i[1817]) | ( l_40 [1417] &  i[1817]);
assign l_39[718]    = ( l_40 [1418] & !i[1817]) | ( l_40 [1419] &  i[1817]);
assign l_39[719]    = ( l_40 [1420] & !i[1817]) | ( l_40 [1421] &  i[1817]);
assign l_39[720]    = ( l_40 [1422] & !i[1817]) | ( l_40 [1423] &  i[1817]);
assign l_39[721]    = ( l_40 [1424] & !i[1817]) | ( l_40 [1425] &  i[1817]);
assign l_39[722]    = ( l_40 [1426] & !i[1817]) | ( l_40 [1427] &  i[1817]);
assign l_39[723]    = ( l_40 [1428] & !i[1817]) | ( l_40 [1429] &  i[1817]);
assign l_39[724]    = ( l_40 [1430] & !i[1817]) | ( l_40 [1431] &  i[1817]);
assign l_39[725]    = ( l_40 [1432] & !i[1817]) | ( l_40 [1433] &  i[1817]);
assign l_39[726]    = ( l_40 [1434] & !i[1817]) | ( l_40 [1435] &  i[1817]);
assign l_39[727]    = ( l_40 [1436] & !i[1817]) | ( l_40 [1437] &  i[1817]);
assign l_39[728]    = ( l_40 [1438] & !i[1817]) | ( l_40 [1439] &  i[1817]);
assign l_39[729]    = ( l_40 [1440] & !i[1817]) | ( l_40 [1441] &  i[1817]);
assign l_39[730]    = ( l_40 [1442] & !i[1817]) | ( l_40 [1443] &  i[1817]);
assign l_39[731]    = ( l_40 [1444] & !i[1817]) | ( l_40 [1445] &  i[1817]);
assign l_39[732]    = ( l_40 [1446] & !i[1817]) | ( l_40 [1447] &  i[1817]);
assign l_39[733]    = ( l_40 [1448] & !i[1817]) | ( l_40 [1449] &  i[1817]);
assign l_39[734]    = ( l_40 [1450] & !i[1817]) | ( l_40 [1451] &  i[1817]);
assign l_39[735]    = ( l_40 [1452] & !i[1817]) | ( l_40 [1453] &  i[1817]);
assign l_39[736]    = ( l_40 [1454] & !i[1817]) | ( l_40 [1455] &  i[1817]);
assign l_39[737]    = ( l_40 [1456] & !i[1817]) | ( l_40 [1457] &  i[1817]);
assign l_39[738]    = ( l_40 [1458] & !i[1817]) | ( l_40 [1459] &  i[1817]);
assign l_39[739]    = ( l_40 [1460] & !i[1817]) | ( l_40 [1461] &  i[1817]);
assign l_39[740]    = ( l_40 [1462] & !i[1817]) | ( l_40 [1463] &  i[1817]);
assign l_39[741]    = ( l_40 [1464] & !i[1817]) | ( l_40 [1465] &  i[1817]);
assign l_39[742]    = ( l_40 [1466] & !i[1817]) | ( l_40 [1467] &  i[1817]);
assign l_39[743]    = ( l_40 [1468] & !i[1817]) | ( l_40 [1469] &  i[1817]);
assign l_39[744]    = ( l_40 [1470] & !i[1817]) | ( l_40 [1471] &  i[1817]);
assign l_39[745]    = ( l_40 [1472] & !i[1817]) | ( l_40 [1473] &  i[1817]);
assign l_39[746]    = ( l_40 [1474] & !i[1817]) | ( l_40 [1475] &  i[1817]);
assign l_39[747]    = ( l_40 [1476] & !i[1817]) | ( l_40 [1477] &  i[1817]);
assign l_39[748]    = ( l_40 [1478] & !i[1817]) | ( l_40 [1479] &  i[1817]);
assign l_39[749]    = ( l_40 [1480] & !i[1817]) | ( l_40 [1481] &  i[1817]);
assign l_39[750]    = ( l_40 [1482] & !i[1817]) | ( l_40 [1483] &  i[1817]);
assign l_39[751]    = ( l_40 [1484] & !i[1817]) | ( l_40 [1485] &  i[1817]);
assign l_39[752]    = ( l_40 [1486] & !i[1817]) | ( l_40 [1487] &  i[1817]);
assign l_39[753]    = ( l_40 [1488] & !i[1817]) | ( l_40 [1489] &  i[1817]);
assign l_39[754]    = ( l_40 [1490] & !i[1817]) | ( l_40 [1491] &  i[1817]);
assign l_39[755]    = ( l_40 [1492] & !i[1817]) | ( l_40 [1493] &  i[1817]);
assign l_39[756]    = ( l_40 [1494] & !i[1817]) | ( l_40 [1495] &  i[1817]);
assign l_39[757]    = ( l_40 [1496] & !i[1817]) | ( l_40 [1497] &  i[1817]);
assign l_39[758]    = ( l_40 [1498] & !i[1817]) | ( l_40 [1499] &  i[1817]);
assign l_39[759]    = ( l_40 [1500] & !i[1817]) | ( l_40 [1501] &  i[1817]);
assign l_39[760]    = ( l_40 [1502] & !i[1817]) | ( l_40 [1503] &  i[1817]);
assign l_39[761]    = ( l_40 [1504] & !i[1817]) | ( l_40 [1505] &  i[1817]);
assign l_39[762]    = ( l_40 [1506] & !i[1817]) | ( l_40 [1507] &  i[1817]);
assign l_39[763]    = ( l_40 [1508] & !i[1817]) | ( l_40 [1509] &  i[1817]);
assign l_39[764]    = ( l_40 [1510] & !i[1817]) | ( l_40 [1511] &  i[1817]);
assign l_39[765]    = ( l_40 [1512] & !i[1817]) | ( l_40 [1513] &  i[1817]);
assign l_39[766]    = ( l_40 [1514] & !i[1817]) | ( l_40 [1515] &  i[1817]);
assign l_39[767]    = ( l_40 [1516] & !i[1817]) | ( l_40 [1517] &  i[1817]);
assign l_39[768]    = ( l_40 [1518] & !i[1817]) | ( l_40 [1519] &  i[1817]);
assign l_39[769]    = ( l_40 [1520] & !i[1817]) | ( l_40 [1521] &  i[1817]);
assign l_39[770]    = ( l_40 [1522] & !i[1817]) | ( l_40 [1523] &  i[1817]);
assign l_39[771]    = ( l_40 [1524] & !i[1817]) | ( l_40 [1525] &  i[1817]);
assign l_39[772]    = ( l_40 [1526] & !i[1817]) | ( l_40 [1527] &  i[1817]);
assign l_39[773]    = ( l_40 [1528] & !i[1817]) | ( l_40 [1529] &  i[1817]);
assign l_39[774]    = ( l_40 [1530] & !i[1817]) | ( l_40 [1531] &  i[1817]);
assign l_39[775]    = ( l_40 [1532] & !i[1817]) | ( l_40 [1533] &  i[1817]);
assign l_39[776]    = ( l_40 [1534] & !i[1817]) | ( l_40 [1535] &  i[1817]);
assign l_39[777]    = ( l_40 [1536] & !i[1817]) | ( l_40 [1537] &  i[1817]);
assign l_39[778]    = ( l_40 [1538] & !i[1817]) | ( l_40 [1539] &  i[1817]);
assign l_39[779]    = ( l_40 [1540] & !i[1817]) | ( l_40 [1541] &  i[1817]);
assign l_39[780]    = ( l_40 [1542] & !i[1817]) | ( l_40 [1543] &  i[1817]);
assign l_39[781]    = ( l_40 [1544] & !i[1817]) | ( l_40 [1545] &  i[1817]);
assign l_39[782]    = ( l_40 [1546] & !i[1817]) | ( l_40 [1547] &  i[1817]);
assign l_39[783]    = ( l_40 [1548] & !i[1817]) | ( l_40 [1549] &  i[1817]);
assign l_39[784]    = ( l_40 [1550] & !i[1817]) | ( l_40 [1551] &  i[1817]);
assign l_39[785]    = ( l_40 [1552] & !i[1817]) | ( l_40 [1553] &  i[1817]);
assign l_39[786]    = ( l_40 [1554] & !i[1817]) | ( l_40 [1555] &  i[1817]);
assign l_39[787]    = ( l_40 [1556] & !i[1817]) | ( l_40 [1557] &  i[1817]);
assign l_39[788]    = ( l_40 [1558] & !i[1817]) | ( l_40 [1559] &  i[1817]);
assign l_39[789]    = ( l_40 [1560] & !i[1817]) | ( l_40 [1561] &  i[1817]);
assign l_39[790]    = ( l_40 [1562] & !i[1817]) | ( l_40 [1563] &  i[1817]);
assign l_39[791]    = ( l_40 [1564] & !i[1817]) | ( l_40 [1565] &  i[1817]);
assign l_39[792]    = ( l_40 [1566] & !i[1817]) | ( l_40 [1567] &  i[1817]);
assign l_39[793]    = ( l_40 [1568] & !i[1817]) | ( l_40 [1569] &  i[1817]);
assign l_39[794]    = ( l_40 [1570] & !i[1817]) | ( l_40 [1571] &  i[1817]);
assign l_39[795]    = ( l_40 [1572] & !i[1817]) | ( l_40 [1573] &  i[1817]);
assign l_39[796]    = ( l_40 [1574] & !i[1817]) | ( l_40 [1575] &  i[1817]);
assign l_39[797]    = ( l_40 [1576] & !i[1817]) | ( l_40 [1577] &  i[1817]);
assign l_39[798]    = ( l_40 [1578] & !i[1817]) | ( l_40 [1579] &  i[1817]);
assign l_39[799]    = ( l_40 [1580] & !i[1817]) | ( l_40 [1581] &  i[1817]);
assign l_39[800]    = ( l_40 [1582] & !i[1817]) | ( l_40 [1583] &  i[1817]);
assign l_39[801]    = ( l_40 [1584] & !i[1817]) | ( l_40 [1585] &  i[1817]);
assign l_39[802]    = ( l_40 [1586] & !i[1817]) | ( l_40 [1587] &  i[1817]);
assign l_39[803]    = ( l_40 [1588] & !i[1817]) | ( l_40 [1589] &  i[1817]);
assign l_39[804]    = ( l_40 [1590] & !i[1817]) | ( l_40 [1591] &  i[1817]);
assign l_39[805]    = ( l_40 [1592] & !i[1817]) | ( l_40 [1593] &  i[1817]);
assign l_39[806]    = ( l_40 [1594] & !i[1817]) | ( l_40 [1595] &  i[1817]);
assign l_39[807]    = ( l_40 [1596] & !i[1817]) | ( l_40 [1597] &  i[1817]);
assign l_39[808]    = ( l_40 [1598] & !i[1817]) | ( l_40 [1599] &  i[1817]);
assign l_39[809]    = ( l_40 [1600] & !i[1817]) | ( l_40 [1601] &  i[1817]);
assign l_39[810]    = ( l_40 [1602] & !i[1817]) | ( l_40 [1603] &  i[1817]);
assign l_39[811]    = ( l_40 [1604] & !i[1817]) | ( l_40 [1605] &  i[1817]);
assign l_39[812]    = ( l_40 [1606] & !i[1817]) | ( l_40 [1607] &  i[1817]);
assign l_39[813]    = ( l_40 [1608] & !i[1817]) | ( l_40 [1609] &  i[1817]);
assign l_39[814]    = ( l_40 [1610] & !i[1817]) | ( l_40 [1611] &  i[1817]);
assign l_39[815]    = ( l_40 [1612] & !i[1817]) | ( l_40 [1613] &  i[1817]);
assign l_39[816]    = ( l_40 [1614] & !i[1817]) | ( l_40 [1615] &  i[1817]);
assign l_39[817]    = ( l_40 [1616] & !i[1817]) | ( l_40 [1617] &  i[1817]);
assign l_39[818]    = ( l_40 [1618] & !i[1817]) | ( l_40 [1619] &  i[1817]);
assign l_39[819]    = ( l_40 [1620] & !i[1817]) | ( l_40 [1621] &  i[1817]);
assign l_39[820]    = ( l_40 [1622] & !i[1817]) | ( l_40 [1623] &  i[1817]);
assign l_39[821]    = ( l_40 [1624] & !i[1817]) | ( l_40 [1625] &  i[1817]);
assign l_39[822]    = ( l_40 [1626] & !i[1817]) | ( l_40 [1627] &  i[1817]);
assign l_39[823]    = ( l_40 [1628] & !i[1817]) | ( l_40 [1629] &  i[1817]);
assign l_39[824]    = ( l_40 [1630] & !i[1817]) | ( l_40 [1631] &  i[1817]);
assign l_39[825]    = ( l_40 [1632] & !i[1817]) | ( l_40 [1633] &  i[1817]);
assign l_39[826]    = ( l_40 [1634] & !i[1817]) | ( l_40 [1635] &  i[1817]);
assign l_39[827]    = ( l_40 [1636] & !i[1817]) | ( l_40 [1637] &  i[1817]);
assign l_39[828]    = ( l_40 [1638] & !i[1817]) | ( l_40 [1639] &  i[1817]);
assign l_39[829]    = ( l_40 [1640] & !i[1817]) | ( l_40 [1641] &  i[1817]);
assign l_39[830]    = ( l_40 [1642] & !i[1817]) | ( l_40 [1643] &  i[1817]);
assign l_39[831]    = ( l_40 [1644] & !i[1817]) | ( l_40 [1645] &  i[1817]);
assign l_39[832]    = ( l_40 [1646] & !i[1817]) | ( l_40 [1647] &  i[1817]);
assign l_39[833]    = ( l_40 [1648] & !i[1817]) | ( l_40 [1649] &  i[1817]);
assign l_39[834]    = ( l_40 [1650] & !i[1817]) | ( l_40 [1651] &  i[1817]);
assign l_39[835]    = ( l_40 [1652] & !i[1817]) | ( l_40 [1653] &  i[1817]);
assign l_39[836]    = ( l_40 [1654] & !i[1817]) | ( l_40 [1655] &  i[1817]);
assign l_39[837]    = ( l_40 [1656] & !i[1817]) | ( l_40 [1657] &  i[1817]);
assign l_39[838]    = ( l_40 [1658] & !i[1817]) | ( l_40 [1659] &  i[1817]);
assign l_39[839]    = ( l_40 [1660] & !i[1817]) | ( l_40 [1661] &  i[1817]);
assign l_39[840]    = ( l_40 [1662] & !i[1817]) | ( l_40 [1663] &  i[1817]);
assign l_39[841]    = ( l_40 [1664] & !i[1817]) | ( l_40 [1665] &  i[1817]);
assign l_39[842]    = ( l_40 [1666] & !i[1817]) | ( l_40 [1667] &  i[1817]);
assign l_39[843]    = ( l_40 [1668] & !i[1817]) | ( l_40 [1669] &  i[1817]);
assign l_39[844]    = ( l_40 [1670] & !i[1817]) | ( l_40 [1671] &  i[1817]);
assign l_39[845]    = ( l_40 [1672] & !i[1817]) | ( l_40 [1673] &  i[1817]);
assign l_39[846]    = ( l_40 [1674] & !i[1817]) | ( l_40 [1675] &  i[1817]);
assign l_39[847]    = ( l_40 [1676] & !i[1817]) | ( l_40 [1677] &  i[1817]);
assign l_39[848]    = ( l_40 [1678] & !i[1817]) | ( l_40 [1679] &  i[1817]);
assign l_39[849]    = ( l_40 [1680] & !i[1817]) | ( l_40 [1681] &  i[1817]);
assign l_39[850]    = ( l_40 [1682] & !i[1817]) | ( l_40 [1683] &  i[1817]);
assign l_39[851]    = ( l_40 [1684] & !i[1817]) | ( l_40 [1685] &  i[1817]);
assign l_39[852]    = ( l_40 [1686] & !i[1817]) | ( l_40 [1687] &  i[1817]);
assign l_39[853]    = ( l_40 [1688] & !i[1817]) | ( l_40 [1689] &  i[1817]);
assign l_39[854]    = ( l_40 [1690] & !i[1817]) | ( l_40 [1691] &  i[1817]);
assign l_39[855]    = ( l_40 [1692] & !i[1817]) | ( l_40 [1693] &  i[1817]);
assign l_39[856]    = ( l_40 [1694] & !i[1817]) | ( l_40 [1695] &  i[1817]);
assign l_39[857]    = ( l_40 [1696] & !i[1817]) | ( l_40 [1697] &  i[1817]);
assign l_39[858]    = ( l_40 [1698] & !i[1817]) | ( l_40 [1699] &  i[1817]);
assign l_39[859]    = ( l_40 [1700] & !i[1817]) | ( l_40 [1701] &  i[1817]);
assign l_39[860]    = ( l_40 [1702] & !i[1817]) | ( l_40 [1703] &  i[1817]);
assign l_39[861]    = ( l_40 [1704] & !i[1817]) | ( l_40 [1705] &  i[1817]);
assign l_39[862]    = ( l_40 [1706] & !i[1817]) | ( l_40 [1707] &  i[1817]);
assign l_39[863]    = ( l_40 [1708] & !i[1817]) | ( l_40 [1709] &  i[1817]);
assign l_39[864]    = ( l_40 [1710] & !i[1817]) | ( l_40 [1711] &  i[1817]);
assign l_39[865]    = ( l_40 [1712] & !i[1817]) | ( l_40 [1713] &  i[1817]);
assign l_39[866]    = ( l_40 [1714] & !i[1817]) | ( l_40 [1715] &  i[1817]);
assign l_39[867]    = ( l_40 [1716] & !i[1817]) | ( l_40 [1717] &  i[1817]);
assign l_39[868]    = ( l_40 [1718] & !i[1817]) | ( l_40 [1719] &  i[1817]);
assign l_39[869]    = ( l_40 [1720] & !i[1817]) | ( l_40 [1721] &  i[1817]);
assign l_39[870]    = ( l_40 [1722] & !i[1817]) | ( l_40 [1723] &  i[1817]);
assign l_39[871]    = ( l_40 [1724] & !i[1817]) | ( l_40 [1725] &  i[1817]);
assign l_39[872]    = ( l_40 [1726] & !i[1817]) | ( l_40 [1727] &  i[1817]);
assign l_39[873]    = ( l_40 [1728] & !i[1817]) | ( l_40 [1729] &  i[1817]);
assign l_39[874]    = ( l_40 [1730] & !i[1817]) | ( l_40 [1731] &  i[1817]);
assign l_39[875]    = ( l_40 [1732] & !i[1817]) | ( l_40 [1733] &  i[1817]);
assign l_39[876]    = ( l_40 [1734] & !i[1817]) | ( l_40 [1735] &  i[1817]);
assign l_39[877]    = ( l_40 [1736] & !i[1817]) | ( l_40 [1737] &  i[1817]);
assign l_39[878]    = ( l_40 [1738] & !i[1817]) | ( l_40 [1739] &  i[1817]);
assign l_39[879]    = ( l_40 [1740] & !i[1817]) | ( l_40 [1741] &  i[1817]);
assign l_39[880]    = ( l_40 [1742] & !i[1817]) | ( l_40 [1743] &  i[1817]);
assign l_39[881]    = ( l_40 [1744] & !i[1817]) | ( l_40 [1745] &  i[1817]);
assign l_39[882]    = ( l_40 [1746] & !i[1817]) | ( l_40 [1747] &  i[1817]);
assign l_39[883]    = ( l_40 [1748] & !i[1817]) | ( l_40 [1749] &  i[1817]);
assign l_39[884]    = ( l_40 [1750] & !i[1817]) | ( l_40 [1751] &  i[1817]);
assign l_39[885]    = ( l_40 [1752] & !i[1817]) | ( l_40 [1753] &  i[1817]);
assign l_39[886]    = ( l_40 [1754] & !i[1817]) | ( l_40 [1755] &  i[1817]);
assign l_39[887]    = ( l_40 [1756] & !i[1817]) | ( l_40 [1757] &  i[1817]);
assign l_39[888]    = ( l_40 [1758] & !i[1817]) | ( l_40 [1759] &  i[1817]);
assign l_39[889]    = ( l_40 [1760] & !i[1817]) | ( l_40 [1761] &  i[1817]);
assign l_39[890]    = ( l_40 [1762] & !i[1817]) | ( l_40 [1763] &  i[1817]);
assign l_39[891]    = ( l_40 [1764] & !i[1817]) | ( l_40 [1765] &  i[1817]);
assign l_39[892]    = ( l_40 [1766] & !i[1817]) | ( l_40 [1767] &  i[1817]);
assign l_39[893]    = ( l_40 [1768] & !i[1817]) | ( l_40 [1769] &  i[1817]);
assign l_39[894]    = ( l_40 [1770] & !i[1817]) | ( l_40 [1771] &  i[1817]);
assign l_39[895]    = ( l_40 [1772] & !i[1817]) | ( l_40 [1773] &  i[1817]);
assign l_39[896]    = ( l_40 [1774] & !i[1817]) | ( l_40 [1775] &  i[1817]);
assign l_39[897]    = ( l_40 [1776] & !i[1817]) | ( l_40 [1777] &  i[1817]);
assign l_39[898]    = ( l_40 [1778] & !i[1817]) | ( l_40 [1779] &  i[1817]);
assign l_39[899]    = ( l_40 [1780] & !i[1817]) | ( l_40 [1781] &  i[1817]);
assign l_39[900]    = ( l_40 [1782] & !i[1817]) | ( l_40 [1783] &  i[1817]);
assign l_39[901]    = ( l_40 [1784] & !i[1817]) | ( l_40 [1785] &  i[1817]);
assign l_39[902]    = ( l_40 [1786] & !i[1817]) | ( l_40 [1787] &  i[1817]);
assign l_39[903]    = ( l_40 [1788] & !i[1817]) | ( l_40 [1789] &  i[1817]);
assign l_39[904]    = ( l_40 [1790] & !i[1817]) | ( l_40 [1791] &  i[1817]);
assign l_39[905]    = ( l_40 [1792] & !i[1817]) | ( l_40 [1793] &  i[1817]);
assign l_39[906]    = ( l_40 [1794] & !i[1817]) | ( l_40 [1795] &  i[1817]);
assign l_39[907]    = ( l_40 [1796] & !i[1817]) | ( l_40 [1797] &  i[1817]);
assign l_39[908]    = ( l_40 [1798] & !i[1817]) | ( l_40 [1799] &  i[1817]);
assign l_39[909]    = ( l_40 [1800] & !i[1817]) | ( l_40 [1801] &  i[1817]);
assign l_39[910]    = ( l_40 [1802] & !i[1817]) | ( l_40 [1803] &  i[1817]);
assign l_39[911]    = ( l_40 [1804] & !i[1817]) | ( l_40 [1805] &  i[1817]);
assign l_39[912]    = ( l_40 [1806] & !i[1817]) | ( l_40 [1807] &  i[1817]);
assign l_39[913]    = ( l_40 [1808] & !i[1817]) | ( l_40 [1809] &  i[1817]);
assign l_39[914]    = ( l_40 [1810] & !i[1817]) | ( l_40 [1811] &  i[1817]);
assign l_39[915]    = ( l_40 [1812] & !i[1817]) | ( l_40 [1813] &  i[1817]);
assign l_39[916]    = ( l_40 [1814] & !i[1817]) | ( l_40 [1815] &  i[1817]);
assign l_39[917]    = ( l_40 [1816] & !i[1817]) | ( l_40 [1817] &  i[1817]);
assign l_39[918]    = ( l_40 [1818] & !i[1817]) | ( l_40 [1819] &  i[1817]);
assign l_39[919]    = ( l_40 [1820] & !i[1817]) | ( l_40 [1821] &  i[1817]);
assign l_39[920]    = ( l_40 [1822] & !i[1817]) | ( l_40 [1823] &  i[1817]);
assign l_39[921]    = ( l_40 [1824] & !i[1817]) | ( l_40 [1825] &  i[1817]);
assign l_39[922]    = ( l_40 [1826] & !i[1817]) | ( l_40 [1827] &  i[1817]);
assign l_39[923]    = ( l_40 [1828] & !i[1817]) | ( l_40 [1829] &  i[1817]);
assign l_39[924]    = ( l_40 [1830] & !i[1817]) | ( l_40 [1831] &  i[1817]);
assign l_39[925]    = ( l_40 [1832] & !i[1817]) | ( l_40 [1833] &  i[1817]);
assign l_39[926]    = ( l_40 [1834] & !i[1817]) | ( l_40 [1835] &  i[1817]);
assign l_39[927]    = ( l_40 [1836] & !i[1817]) | ( l_40 [1837] &  i[1817]);
assign l_39[928]    = ( l_40 [1838] & !i[1817]) | ( l_40 [1839] &  i[1817]);
assign l_39[929]    = ( l_40 [1840] & !i[1817]) | ( l_40 [1841] &  i[1817]);
assign l_39[930]    = ( l_40 [1842] & !i[1817]) | ( l_40 [1843] &  i[1817]);
assign l_39[931]    = ( l_40 [1844] & !i[1817]) | ( l_40 [1845] &  i[1817]);
assign l_39[932]    = ( l_40 [1846] & !i[1817]) | ( l_40 [1847] &  i[1817]);
assign l_39[933]    = ( l_40 [1848] & !i[1817]) | ( l_40 [1849] &  i[1817]);
assign l_39[934]    = ( l_40 [1850] & !i[1817]) | ( l_40 [1851] &  i[1817]);
assign l_39[935]    = ( l_40 [1852] & !i[1817]) | ( l_40 [1853] &  i[1817]);
assign l_39[936]    = ( l_40 [1854] & !i[1817]) | ( l_40 [1855] &  i[1817]);
assign l_39[937]    = ( l_40 [1856] & !i[1817]) | ( l_40 [1857] &  i[1817]);
assign l_39[938]    = ( l_40 [1858] & !i[1817]) | ( l_40 [1859] &  i[1817]);
assign l_39[939]    = ( l_40 [1860] & !i[1817]) | ( l_40 [1861] &  i[1817]);
assign l_39[940]    = ( l_40 [1862] & !i[1817]) | ( l_40 [1863] &  i[1817]);
assign l_39[941]    = ( l_40 [1864] & !i[1817]) | ( l_40 [1865] &  i[1817]);
assign l_39[942]    = ( l_40 [1866] & !i[1817]) | ( l_40 [1867] &  i[1817]);
assign l_39[943]    = ( l_40 [1868] & !i[1817]) | ( l_40 [1869] &  i[1817]);
assign l_39[944]    = ( l_40 [1870] & !i[1817]) | ( l_40 [1871] &  i[1817]);
assign l_39[945]    = ( l_40 [1872] & !i[1817]) | ( l_40 [1873] &  i[1817]);
assign l_39[946]    = ( l_40 [1874] & !i[1817]) | ( l_40 [1875] &  i[1817]);
assign l_39[947]    = ( l_40 [1876] & !i[1817]) | ( l_40 [1877] &  i[1817]);
assign l_39[948]    = ( l_40 [1878] & !i[1817]) | ( l_40 [1879] &  i[1817]);
assign l_39[949]    = ( l_40 [1880] & !i[1817]) | ( l_40 [1881] &  i[1817]);
assign l_39[950]    = ( l_40 [1882] & !i[1817]) | ( l_40 [1883] &  i[1817]);
assign l_39[951]    = ( l_40 [1884] & !i[1817]) | ( l_40 [1885] &  i[1817]);
assign l_39[952]    = ( l_40 [1886] & !i[1817]) | ( l_40 [1887] &  i[1817]);
assign l_39[953]    = ( l_40 [1888] & !i[1817]) | ( l_40 [1889] &  i[1817]);
assign l_39[954]    = ( l_40 [1890] & !i[1817]) | ( l_40 [1891] &  i[1817]);
assign l_39[955]    = ( l_40 [1892] & !i[1817]) | ( l_40 [1893] &  i[1817]);
assign l_39[956]    = ( l_40 [1894] & !i[1817]) | ( l_40 [1895] &  i[1817]);
assign l_39[957]    = ( l_40 [1896] & !i[1817]) | ( l_40 [1897] &  i[1817]);
assign l_39[958]    = ( l_40 [1898] & !i[1817]) | ( l_40 [1899] &  i[1817]);
assign l_39[959]    = ( l_40 [1900] & !i[1817]) | ( l_40 [1901] &  i[1817]);
assign l_39[960]    = ( l_40 [1902] & !i[1817]) | ( l_40 [1903] &  i[1817]);
assign l_39[961]    = ( l_40 [1904] & !i[1817]) | ( l_40 [1905] &  i[1817]);
assign l_39[962]    = ( l_40 [1906] & !i[1817]) | ( l_40 [1907] &  i[1817]);
assign l_39[963]    = ( l_40 [1908] & !i[1817]) | ( l_40 [1909] &  i[1817]);
assign l_39[964]    = ( l_40 [1910] & !i[1817]) | ( l_40 [1911] &  i[1817]);
assign l_39[965]    = ( l_40 [1912] & !i[1817]) | ( l_40 [1913] &  i[1817]);
assign l_39[966]    = ( l_40 [1914] & !i[1817]) | ( l_40 [1915] &  i[1817]);
assign l_39[967]    = ( l_40 [1916] & !i[1817]) | ( l_40 [1917] &  i[1817]);
assign l_39[968]    = ( l_40 [1918] & !i[1817]) | ( l_40 [1919] &  i[1817]);
assign l_39[969]    = ( l_40 [1920] & !i[1817]) | ( l_40 [1921] &  i[1817]);
assign l_39[970]    = ( l_40 [1922] & !i[1817]) | ( l_40 [1923] &  i[1817]);
assign l_39[971]    = ( l_40 [1924] & !i[1817]) | ( l_40 [1925] &  i[1817]);
assign l_39[972]    = ( l_40 [1926] & !i[1817]) | ( l_40 [1927] &  i[1817]);
assign l_39[973]    = ( l_40 [1928] & !i[1817]) | ( l_40 [1929] &  i[1817]);
assign l_39[974]    = ( l_40 [1930] & !i[1817]) | ( l_40 [1931] &  i[1817]);
assign l_39[975]    = ( l_40 [1932] & !i[1817]) | ( l_40 [1933] &  i[1817]);
assign l_39[976]    = ( l_40 [1934] & !i[1817]) | ( l_40 [1935] &  i[1817]);
assign l_39[977]    = ( l_40 [1936] & !i[1817]) | ( l_40 [1937] &  i[1817]);
assign l_39[978]    = ( l_40 [1938] & !i[1817]) | ( l_40 [1939] &  i[1817]);
assign l_39[979]    = ( l_40 [1940] & !i[1817]) | ( l_40 [1941] &  i[1817]);
assign l_39[980]    = ( l_40 [1942] & !i[1817]) | ( l_40 [1943] &  i[1817]);
assign l_39[981]    = ( l_40 [1944] & !i[1817]) | ( l_40 [1945] &  i[1817]);
assign l_39[982]    = ( l_40 [1946] & !i[1817]) | ( l_40 [1947] &  i[1817]);
assign l_39[983]    = ( l_40 [1948] & !i[1817]) | ( l_40 [1949] &  i[1817]);
assign l_39[984]    = ( l_40 [1950] & !i[1817]) | ( l_40 [1951] &  i[1817]);
assign l_39[985]    = ( l_40 [1952] & !i[1817]) | ( l_40 [1953] &  i[1817]);
assign l_39[986]    = ( l_40 [1954] & !i[1817]) | ( l_40 [1955] &  i[1817]);
assign l_39[987]    = ( l_40 [1956] & !i[1817]) | ( l_40 [1957] &  i[1817]);
assign l_39[988]    = ( l_40 [1958] & !i[1817]) | ( l_40 [1959] &  i[1817]);
assign l_39[989]    = ( l_40 [1960] & !i[1817]) | ( l_40 [1961] &  i[1817]);
assign l_39[990]    = ( l_40 [1962] & !i[1817]) | ( l_40 [1963] &  i[1817]);
assign l_39[991]    = ( l_40 [1964] & !i[1817]) | ( l_40 [1965] &  i[1817]);
assign l_39[992]    = ( l_40 [1966] & !i[1817]) | ( l_40 [1967] &  i[1817]);
assign l_39[993]    = ( l_40 [1968] & !i[1817]) | ( l_40 [1969] &  i[1817]);
assign l_39[994]    = ( l_40 [1970] & !i[1817]) | ( l_40 [1971] &  i[1817]);
assign l_39[995]    = ( l_40 [1972] & !i[1817]) | ( l_40 [1973] &  i[1817]);
assign l_39[996]    = ( l_40 [1974] & !i[1817]) | ( l_40 [1975] &  i[1817]);
assign l_39[997]    = ( l_40 [1976] & !i[1817]) | ( l_40 [1977] &  i[1817]);
assign l_39[998]    = ( l_40 [1978] & !i[1817]) | ( l_40 [1979] &  i[1817]);
assign l_39[999]    = ( l_40 [1980] & !i[1817]) | ( l_40 [1981] &  i[1817]);
assign l_39[1000]    = ( l_40 [1982] & !i[1817]) | ( l_40 [1983] &  i[1817]);
assign l_39[1001]    = ( l_40 [1984] & !i[1817]) | ( l_40 [1985] &  i[1817]);
assign l_39[1002]    = ( l_40 [1986] & !i[1817]) | ( l_40 [1987] &  i[1817]);
assign l_39[1003]    = ( l_40 [1988] & !i[1817]) | ( l_40 [1989] &  i[1817]);
assign l_39[1004]    = ( l_40 [1990] & !i[1817]) | ( l_40 [1991] &  i[1817]);
assign l_39[1005]    = ( l_40 [1992] & !i[1817]) | ( l_40 [1993] &  i[1817]);
assign l_39[1006]    = ( l_40 [1994] & !i[1817]) | ( l_40 [1995] &  i[1817]);
assign l_39[1007]    = ( l_40 [1996] & !i[1817]) | ( l_40 [1997] &  i[1817]);
assign l_39[1008]    = ( l_40 [1998] & !i[1817]) | ( l_40 [1999] &  i[1817]);
assign l_39[1009]    = ( l_40 [2000] & !i[1817]) | ( l_40 [2001] &  i[1817]);
assign l_39[1010]    = ( l_40 [2002] & !i[1817]) | ( l_40 [2003] &  i[1817]);
assign l_39[1011]    = ( l_40 [2004] & !i[1817]) | ( l_40 [2005] &  i[1817]);
assign l_39[1012]    = ( l_40 [2006] & !i[1817]) | ( l_40 [2007] &  i[1817]);
assign l_39[1013]    = ( l_40 [2008] & !i[1817]) | ( l_40 [2009] &  i[1817]);
assign l_39[1014]    = ( l_40 [2010] & !i[1817]) | ( l_40 [2011] &  i[1817]);
assign l_39[1015]    = ( l_40 [2012] & !i[1817]) | ( l_40 [2013] &  i[1817]);
assign l_39[1016]    = ( l_40 [2014] & !i[1817]) | ( l_40 [2015] &  i[1817]);
assign l_39[1017]    = ( l_40 [2016] & !i[1817]) | ( l_40 [2017] &  i[1817]);
assign l_39[1018]    = ( l_40 [2018] & !i[1817]) | ( l_40 [2019] &  i[1817]);
assign l_39[1019]    = ( l_40 [2020] & !i[1817]) | ( l_40 [2021] &  i[1817]);
assign l_39[1020]    = ( l_40 [2022] & !i[1817]) | ( l_40 [2023] &  i[1817]);
assign l_39[1021]    = ( l_40 [2024] & !i[1817]) | ( l_40 [2025] &  i[1817]);
assign l_39[1022]    = ( l_40 [2026] & !i[1817]) | ( l_40 [2027] &  i[1817]);
assign l_39[1023]    = ( l_40 [2028] & !i[1817]) | ( l_40 [2029] &  i[1817]);
assign l_39[1024]    = ( l_40 [2030] & !i[1817]) | ( l_40 [2031] &  i[1817]);
assign l_39[1025]    = ( l_40 [2032] & !i[1817]) | ( l_40 [2033] &  i[1817]);
assign l_39[1026]    = ( l_40 [2034] & !i[1817]) | ( l_40 [2035] &  i[1817]);
assign l_39[1027]    = ( l_40 [2036] & !i[1817]) | ( l_40 [2037] &  i[1817]);
assign l_39[1028]    = ( l_40 [2038] & !i[1817]) | ( l_40 [2039] &  i[1817]);
assign l_39[1029]    = ( l_40 [2040] & !i[1817]) | ( l_40 [2041] &  i[1817]);
assign l_39[1030]    = ( l_40 [2042] & !i[1817]) | ( l_40 [2043] &  i[1817]);
assign l_39[1031]    = ( l_40 [2044] & !i[1817]) | ( l_40 [2045] &  i[1817]);
assign l_39[1032]    = ( l_40 [2046] & !i[1817]) | ( l_40 [2047] &  i[1817]);
assign l_39[1033]    = ( l_40 [2048] & !i[1817]) | ( l_40 [2049] &  i[1817]);
assign l_39[1034]    = ( l_40 [2050] & !i[1817]) | ( l_40 [2051] &  i[1817]);
assign l_39[1035]    = ( l_40 [2052] & !i[1817]) | ( l_40 [2053] &  i[1817]);
assign l_39[1036]    = ( l_40 [2054] & !i[1817]) | ( l_40 [2055] &  i[1817]);
assign l_39[1037]    = ( l_40 [2056] & !i[1817]) | ( l_40 [2057] &  i[1817]);
assign l_39[1038]    = ( l_40 [2058] & !i[1817]) | ( l_40 [2059] &  i[1817]);
assign l_39[1039]    = ( l_40 [2060] & !i[1817]) | ( l_40 [2061] &  i[1817]);
assign l_39[1040]    = ( l_40 [2062] & !i[1817]) | ( l_40 [2063] &  i[1817]);
assign l_39[1041]    = ( l_40 [2064] & !i[1817]) | ( l_40 [2065] &  i[1817]);
assign l_39[1042]    = ( l_40 [2066]);
assign l_39[1043]    = ( l_40 [2067]);
assign l_39[1044]    = ( l_40 [2068]);
assign l_39[1045]    = ( l_40 [2069]);
assign l_39[1046]    = ( l_40 [2070]);
assign l_39[1047]    = ( l_40 [2071]);
assign l_39[1048]    = ( l_40 [2072]);
assign l_39[1049]    = ( l_40 [2073]);
assign l_39[1050]    = ( l_40 [2074]);
assign l_39[1051]    = ( l_40 [2075]);
assign l_39[1052]    = ( l_40 [2076]);
assign l_39[1053]    = ( l_40 [2077]);
assign l_39[1054]    = ( l_40 [2078]);
assign l_39[1055]    = ( l_40 [2079]);
assign l_39[1056]    = ( l_40 [2080]);
assign l_39[1057]    = ( l_40 [2081]);
assign l_39[1058]    = ( l_40 [2082]);
assign l_39[1059]    = ( l_40 [2083]);
assign l_39[1060]    = ( l_40 [2084]);
assign l_39[1061]    = ( l_40 [2085]);
assign l_39[1062]    = ( l_40 [2086]);
assign l_39[1063]    = ( l_40 [2087]);
assign l_39[1064]    = ( l_40 [2088]);
assign l_39[1065]    = ( l_40 [2089]);
assign l_39[1066]    = ( l_40 [2090]);
assign l_39[1067]    = ( l_40 [2091]);
assign l_39[1068]    = ( l_40 [2092]);
assign l_39[1069]    = ( l_40 [2093]);
assign l_39[1070]    = ( l_40 [2094]);
assign l_39[1071]    = ( l_40 [2095]);
assign l_39[1072]    = ( l_40 [2096]);
assign l_39[1073]    = ( l_40 [2097]);
assign l_39[1074]    = ( l_40 [2098]);
assign l_39[1075]    = ( l_40 [2099]);
assign l_39[1076]    = ( l_40 [2100]);
assign l_39[1077]    = ( l_40 [2101]);
assign l_39[1078]    = ( l_40 [2102]);
assign l_39[1079]    = ( l_40 [2103]);
assign l_39[1080]    = ( l_40 [2104]);
assign l_39[1081]    = ( l_40 [2105]);
assign l_39[1082]    = ( l_40 [2106]);
assign l_39[1083]    = ( l_40 [2107]);
assign l_39[1084]    = ( l_40 [2108]);
assign l_39[1085]    = ( l_40 [2109]);
assign l_39[1086]    = ( l_40 [2110]);
assign l_39[1087]    = ( l_40 [2111]);
assign l_39[1088]    = ( l_40 [2112]);
assign l_39[1089]    = ( l_40 [2113]);
assign l_39[1090]    = ( l_40 [2114]);
assign l_39[1091]    = ( l_40 [2115]);
assign l_39[1092]    = ( l_40 [2116]);
assign l_39[1093]    = ( l_40 [2117]);
assign l_39[1094]    = ( l_40 [2118]);
assign l_39[1095]    = ( l_40 [2119]);
assign l_39[1096]    = ( l_40 [2120]);
assign l_39[1097]    = ( l_40 [2121]);
assign l_39[1098]    = ( l_40 [2122]);
assign l_39[1099]    = ( l_40 [2123]);
assign l_39[1100]    = ( l_40 [2124]);
assign l_39[1101]    = ( l_40 [2125]);
assign l_39[1102]    = ( l_40 [2126]);
assign l_39[1103]    = ( l_40 [2127]);
assign l_39[1104]    = ( l_40 [2128]);
assign l_39[1105]    = ( l_40 [2129]);
assign l_39[1106]    = ( l_40 [2130]);
assign l_39[1107]    = ( l_40 [2131]);
assign l_39[1108]    = ( l_40 [2132]);
assign l_39[1109]    = ( l_40 [2133]);
assign l_39[1110]    = ( l_40 [2134]);
assign l_39[1111]    = ( l_40 [2135]);
assign l_39[1112]    = ( l_40 [2136]);
assign l_39[1113]    = ( l_40 [2137]);
assign l_39[1114]    = ( l_40 [2138]);
assign l_39[1115]    = ( l_40 [2139]);
assign l_39[1116]    = ( l_40 [2140]);
assign l_39[1117]    = ( l_40 [2141]);
assign l_39[1118]    = ( l_40 [2142]);
assign l_39[1119]    = ( l_40 [2143]);
assign l_39[1120]    = ( l_40 [2144]);
assign l_39[1121]    = ( l_40 [2145]);
assign l_39[1122]    = ( l_40 [2146]);
assign l_39[1123]    = ( l_40 [2147]);
assign l_39[1124]    = ( l_40 [2148]);
assign l_39[1125]    = ( l_40 [2149]);
assign l_39[1126]    = ( l_40 [2150]);
assign l_39[1127]    = ( l_40 [2151]);
assign l_39[1128]    = ( l_40 [2152]);
assign l_39[1129]    = ( l_40 [2153]);
assign l_39[1130]    = ( l_40 [2154]);
assign l_39[1131]    = ( l_40 [2155]);
assign l_39[1132]    = ( l_40 [2156]);
assign l_39[1133]    = ( l_40 [2157]);
assign l_39[1134]    = ( l_40 [2158]);
assign l_39[1135]    = ( l_40 [2159]);
assign l_39[1136]    = ( l_40 [2160]);
assign l_39[1137]    = ( l_40 [2161]);
assign l_39[1138]    = ( l_40 [2162]);
assign l_39[1139]    = ( l_40 [2163]);
assign l_39[1140]    = ( l_40 [2164]);
assign l_39[1141]    = ( l_40 [2165]);
assign l_39[1142]    = ( l_40 [2166]);
assign l_39[1143]    = ( l_40 [2167]);
assign l_39[1144]    = ( l_40 [2168]);
assign l_39[1145]    = ( l_40 [2169]);
assign l_39[1146]    = ( l_40 [2170]);
assign l_39[1147]    = ( l_40 [2171]);
assign l_39[1148]    = ( l_40 [2172]);
assign l_39[1149]    = ( l_40 [2173]);
assign l_39[1150]    = ( l_40 [2174]);
assign l_39[1151]    = ( l_40 [2175]);
assign l_39[1152]    = ( l_40 [2176]);
assign l_39[1153]    = ( l_40 [2177]);
assign l_39[1154]    = ( l_40 [2178]);
assign l_39[1155]    = ( l_40 [2179]);
assign l_39[1156]    = ( l_40 [2180]);
assign l_39[1157]    = ( l_40 [2181]);
assign l_39[1158]    = ( l_40 [2182]);
assign l_39[1159]    = ( l_40 [2183]);
assign l_39[1160]    = ( l_40 [2184]);
assign l_39[1161]    = ( l_40 [2185]);
assign l_39[1162]    = ( l_40 [2186]);
assign l_39[1163]    = ( l_40 [2187]);
assign l_39[1164]    = ( l_40 [2188]);
assign l_39[1165]    = ( l_40 [2189]);
assign l_39[1166]    = ( l_40 [2190]);
assign l_39[1167]    = ( l_40 [2191]);
assign l_39[1168]    = ( l_40 [2192]);
assign l_39[1169]    = ( l_40 [2193]);
assign l_39[1170]    = ( l_40 [2194]);
assign l_39[1171]    = ( l_40 [2195]);
assign l_39[1172]    = ( l_40 [2196]);
assign l_39[1173]    = ( l_40 [2197]);
assign l_39[1174]    = ( l_40 [2198]);
assign l_39[1175]    = ( l_40 [2199]);
assign l_39[1176]    = ( l_40 [2200]);
assign l_39[1177]    = ( l_40 [2201]);
assign l_39[1178]    = ( l_40 [2202]);
assign l_39[1179]    = ( l_40 [2203]);
assign l_39[1180]    = ( l_40 [2204]);
assign l_39[1181]    = ( l_40 [2205]);
assign l_39[1182]    = ( l_40 [2206]);
assign l_39[1183]    = ( l_40 [2207]);
assign l_39[1184]    = ( l_40 [2208]);
assign l_39[1185]    = ( l_40 [2209]);
assign l_39[1186]    = ( l_40 [2210]);
assign l_39[1187]    = ( l_40 [2211]);
assign l_39[1188]    = ( l_40 [2212]);
assign l_39[1189]    = ( l_40 [2213]);
assign l_39[1190]    = ( l_40 [2214]);
assign l_39[1191]    = ( l_40 [2215]);
assign l_39[1192]    = ( l_40 [2216]);
assign l_39[1193]    = ( l_40 [2217]);
assign l_39[1194]    = ( l_40 [2218]);
assign l_39[1195]    = ( l_40 [2219]);
assign l_39[1196]    = ( l_40 [2220]);
assign l_39[1197]    = ( l_40 [2221]);
assign l_39[1198]    = ( l_40 [2222]);
assign l_39[1199]    = ( l_40 [2223]);
assign l_39[1200]    = ( l_40 [2224]);
assign l_39[1201]    = ( l_40 [2225]);
assign l_39[1202]    = ( l_40 [2226]);
assign l_39[1203]    = ( l_40 [2227]);
assign l_39[1204]    = ( l_40 [2228]);
assign l_39[1205]    = ( l_40 [2229]);
assign l_39[1206]    = ( l_40 [2230]);
assign l_39[1207]    = ( l_40 [2231]);
assign l_39[1208]    = ( l_40 [2232]);
assign l_39[1209]    = ( l_40 [2233]);
assign l_39[1210]    = ( l_40 [2234]);
assign l_39[1211]    = ( l_40 [2235]);
assign l_39[1212]    = ( l_40 [2236]);
assign l_39[1213]    = ( l_40 [2237]);
assign l_39[1214]    = ( l_40 [2238]);
assign l_39[1215]    = ( l_40 [2239]);
assign l_39[1216]    = ( l_40 [2240]);
assign l_39[1217]    = ( l_40 [2241]);
assign l_39[1218]    = ( l_40 [2242]);
assign l_39[1219]    = ( l_40 [2243]);
assign l_39[1220]    = ( l_40 [2244]);
assign l_39[1221]    = ( l_40 [2245]);
assign l_39[1222]    = ( l_40 [2246]);
assign l_39[1223]    = ( l_40 [2247]);
assign l_39[1224]    = ( l_40 [2248]);
assign l_39[1225]    = ( l_40 [2249]);
assign l_39[1226]    = ( l_40 [2250]);
assign l_39[1227]    = ( l_40 [2251]);
assign l_39[1228]    = ( l_40 [2252]);
assign l_39[1229]    = ( l_40 [2253]);
assign l_39[1230]    = ( l_40 [2254]);
assign l_39[1231]    = ( l_40 [2255]);
assign l_39[1232]    = ( l_40 [2256]);
assign l_39[1233]    = ( l_40 [2257]);
assign l_39[1234]    = ( l_40 [2258]);
assign l_39[1235]    = ( l_40 [2259]);
assign l_39[1236]    = ( l_40 [2260]);
assign l_39[1237]    = ( l_40 [2261]);
assign l_39[1238]    = ( l_40 [2262]);
assign l_39[1239]    = ( l_40 [2263]);
assign l_39[1240]    = ( l_40 [2264]);
assign l_39[1241]    = ( l_40 [2265]);
assign l_39[1242]    = ( l_40 [2266]);
assign l_39[1243]    = ( l_40 [2267]);
assign l_39[1244]    = ( l_40 [2268]);
assign l_39[1245]    = ( l_40 [2269]);
assign l_39[1246]    = ( l_40 [2270]);
assign l_39[1247]    = ( l_40 [2271]);
assign l_39[1248]    = ( l_40 [2272]);
assign l_39[1249]    = ( l_40 [2273]);
assign l_39[1250]    = ( l_40 [2274]);
assign l_39[1251]    = ( l_40 [2275]);
assign l_39[1252]    = ( l_40 [2276]);
assign l_39[1253]    = ( l_40 [2277]);
assign l_39[1254]    = ( l_40 [2278]);
assign l_39[1255]    = ( l_40 [2279]);
assign l_39[1256]    = ( l_40 [2280]);
assign l_39[1257]    = ( l_40 [2281]);
assign l_39[1258]    = ( l_40 [2282]);
assign l_39[1259]    = ( l_40 [2283]);
assign l_39[1260]    = ( l_40 [2284]);
assign l_39[1261]    = ( l_40 [2285]);
assign l_39[1262]    = ( l_40 [2286]);
assign l_39[1263]    = ( l_40 [2287]);
assign l_39[1264]    = ( l_40 [2288]);
assign l_39[1265]    = ( l_40 [2289]);
assign l_39[1266]    = ( l_40 [2290]);
assign l_39[1267]    = ( l_40 [2291]);
assign l_39[1268]    = ( l_40 [2292]);
assign l_39[1269]    = ( l_40 [2293]);
assign l_39[1270]    = ( l_40 [2294]);
assign l_39[1271]    = ( l_40 [2295]);
assign l_39[1272]    = ( l_40 [2296]);
assign l_39[1273]    = ( l_40 [2297]);
assign l_39[1274]    = ( l_40 [2298]);
assign l_39[1275]    = ( l_40 [2299]);
assign l_39[1276]    = ( l_40 [2300]);
assign l_39[1277]    = ( l_40 [2301]);
assign l_39[1278]    = ( l_40 [2302]);
assign l_39[1279]    = ( l_40 [2303]);
assign l_39[1280]    = ( l_40 [2304]);
assign l_39[1281]    = ( l_40 [2305]);
assign l_39[1282]    = ( l_40 [2306]);
assign l_39[1283]    = ( l_40 [2307]);
assign l_39[1284]    = ( l_40 [2308]);
assign l_39[1285]    = ( l_40 [2309]);
assign l_39[1286]    = ( l_40 [2310]);
assign l_39[1287]    = ( l_40 [2311]);
assign l_39[1288]    = ( l_40 [2312]);
assign l_39[1289]    = ( l_40 [2313]);
assign l_39[1290]    = ( l_40 [2314]);
assign l_39[1291]    = ( l_40 [2315]);
assign l_39[1292]    = ( l_40 [2316]);
assign l_39[1293]    = ( l_40 [2317]);
assign l_39[1294]    = ( l_40 [2318]);
assign l_39[1295]    = ( l_40 [2319]);
assign l_39[1296]    = ( l_40 [2320]);
assign l_39[1297]    = ( l_40 [2321]);
assign l_39[1298]    = ( l_40 [2322]);
assign l_39[1299]    = ( l_40 [2323]);
assign l_39[1300]    = ( l_40 [2324]);
assign l_39[1301]    = ( l_40 [2325]);
assign l_39[1302]    = ( l_40 [2326]);
assign l_39[1303]    = ( l_40 [2327]);
assign l_39[1304]    = ( l_40 [2328]);
assign l_39[1305]    = ( l_40 [2329]);
assign l_39[1306]    = ( l_40 [2330]);
assign l_39[1307]    = ( l_40 [2331]);
assign l_39[1308]    = ( l_40 [2332]);
assign l_39[1309]    = ( l_40 [2333]);
assign l_39[1310]    = ( l_40 [2334]);
assign l_39[1311]    = ( l_40 [2335]);
assign l_39[1312]    = ( l_40 [2336]);
assign l_39[1313]    = ( l_40 [2337]);
assign l_39[1314]    = ( l_40 [2338]);
assign l_39[1315]    = ( l_40 [2339]);
assign l_39[1316]    = ( l_40 [2340]);
assign l_39[1317]    = ( l_40 [2341]);
assign l_39[1318]    = ( l_40 [2342]);
assign l_39[1319]    = ( l_40 [2343]);
assign l_39[1320]    = ( l_40 [2344]);
assign l_39[1321]    = ( l_40 [2345]);
assign l_39[1322]    = ( l_40 [2346]);
assign l_39[1323]    = ( l_40 [2347]);
assign l_39[1324]    = ( l_40 [2348]);
assign l_39[1325]    = ( l_40 [2349]);
assign l_39[1326]    = ( l_40 [2350]);
assign l_39[1327]    = ( l_40 [2351]);
assign l_39[1328]    = ( l_40 [2352]);
assign l_39[1329]    = ( l_40 [2353]);
assign l_39[1330]    = ( l_40 [2354]);
assign l_39[1331]    = ( l_40 [2355]);
assign l_39[1332]    = ( l_40 [2356]);
assign l_39[1333]    = ( l_40 [2357]);
assign l_39[1334]    = ( l_40 [2358]);
assign l_39[1335]    = ( l_40 [2359]);
assign l_39[1336]    = ( l_40 [2360]);
assign l_39[1337]    = ( l_40 [2361]);
assign l_39[1338]    = ( l_40 [2362]);
assign l_39[1339]    = ( l_40 [2363]);
assign l_39[1340]    = ( l_40 [2364]);
assign l_39[1341]    = ( l_40 [2365]);
assign l_39[1342]    = ( l_40 [2366]);
assign l_39[1343]    = ( l_40 [2367]);
assign l_39[1344]    = ( l_40 [2368]);
assign l_39[1345]    = ( l_40 [2369]);
assign l_39[1346]    = ( l_40 [2370]);
assign l_39[1347]    = ( l_40 [2371]);
assign l_39[1348]    = ( l_40 [2372]);
assign l_39[1349]    = ( l_40 [2373]);
assign l_39[1350]    = ( l_40 [2374]);
assign l_39[1351]    = ( l_40 [2375]);
assign l_39[1352]    = ( l_40 [2376]);
assign l_39[1353]    = ( l_40 [2377]);
assign l_39[1354]    = ( l_40 [2378]);
assign l_39[1355]    = ( l_40 [2379]);
assign l_39[1356]    = ( l_40 [2380]);
assign l_39[1357]    = ( l_40 [2381]);
assign l_39[1358]    = ( l_40 [2382]);
assign l_39[1359]    = ( l_40 [2383]);
assign l_39[1360]    = ( l_40 [2384]);
assign l_39[1361]    = ( l_40 [2385]);
assign l_39[1362]    = ( l_40 [2386]);
assign l_39[1363]    = ( l_40 [2387]);
assign l_39[1364]    = ( l_40 [2388]);
assign l_39[1365]    = ( l_40 [2389]);
assign l_39[1366]    = ( l_40 [2390]);
assign l_39[1367]    = ( l_40 [2391]);
assign l_39[1368]    = ( l_40 [2392]);
assign l_39[1369]    = ( l_40 [2393]);
assign l_39[1370]    = ( l_40 [2394]);
assign l_39[1371]    = ( l_40 [2395]);
assign l_39[1372]    = ( l_40 [2396]);
assign l_39[1373]    = ( l_40 [2397]);
assign l_39[1374]    = ( l_40 [2398]);
assign l_39[1375]    = ( l_40 [2399]);
assign l_39[1376]    = ( l_40 [2400]);
assign l_39[1377]    = ( l_40 [2401]);
assign l_39[1378]    = ( l_40 [2402]);
assign l_39[1379]    = ( l_40 [2403]);
assign l_39[1380]    = ( l_40 [2404]);
assign l_39[1381]    = ( l_40 [2405]);
assign l_39[1382]    = ( l_40 [2406]);
assign l_39[1383]    = ( l_40 [2407]);
assign l_39[1384]    = ( l_40 [2408]);
assign l_39[1385]    = ( l_40 [2409]);
assign l_39[1386]    = ( l_40 [2410]);
assign l_39[1387]    = ( l_40 [2411]);
assign l_39[1388]    = ( l_40 [2412]);
assign l_39[1389]    = ( l_40 [2413]);
assign l_39[1390]    = ( l_40 [2414]);
assign l_39[1391]    = ( l_40 [2415]);
assign l_39[1392]    = ( l_40 [2416]);
assign l_39[1393]    = ( l_40 [2417]);
assign l_39[1394]    = ( l_40 [2418]);
assign l_39[1395]    = ( l_40 [2419]);
assign l_39[1396]    = ( l_40 [2420]);
assign l_39[1397]    = ( l_40 [2421]);
assign l_39[1398]    = ( l_40 [2422]);
assign l_39[1399]    = ( l_40 [2423]);
assign l_39[1400]    = ( l_40 [2424]);
assign l_39[1401]    = ( l_40 [2425]);
assign l_39[1402]    = ( l_40 [2426]);
assign l_39[1403]    = ( l_40 [2427]);
assign l_39[1404]    = ( l_40 [2428]);
assign l_39[1405]    = ( l_40 [2429]);
assign l_39[1406]    = ( l_40 [2430]);
assign l_39[1407]    = ( l_40 [2431]);
assign l_39[1408]    = ( l_40 [2432]);
assign l_39[1409]    = ( l_40 [2433]);
assign l_39[1410]    = ( l_40 [2434]);
assign l_39[1411]    = ( l_40 [2435]);
assign l_39[1412]    = ( l_40 [2436]);
assign l_39[1413]    = ( l_40 [2437]);
assign l_39[1414]    = ( l_40 [2438]);
assign l_39[1415]    = ( l_40 [2439]);
assign l_39[1416]    = ( l_40 [2440]);
assign l_39[1417]    = ( l_40 [2441]);
assign l_39[1418]    = ( l_40 [2442]);
assign l_39[1419]    = ( l_40 [2443]);
assign l_39[1420]    = ( l_40 [2444]);
assign l_39[1421]    = ( l_40 [2445]);
assign l_39[1422]    = ( l_40 [2446]);
assign l_39[1423]    = ( l_40 [2447]);
assign l_39[1424]    = ( l_40 [2448]);
assign l_39[1425]    = ( l_40 [2449]);
assign l_39[1426]    = ( l_40 [2450]);
assign l_39[1427]    = ( l_40 [2451]);
assign l_39[1428]    = ( l_40 [2452]);
assign l_39[1429]    = ( l_40 [2453]);
assign l_39[1430]    = ( l_40 [2454]);
assign l_39[1431]    = ( l_40 [2455]);
assign l_39[1432]    = ( l_40 [2456]);
assign l_39[1433]    = ( l_40 [2457]);
assign l_39[1434]    = ( l_40 [2458]);
assign l_39[1435]    = ( l_40 [2459]);
assign l_39[1436]    = ( l_40 [2460]);
assign l_39[1437]    = ( l_40 [2461]);
assign l_39[1438]    = ( l_40 [2462]);
assign l_39[1439]    = ( l_40 [2463]);
assign l_39[1440]    = ( l_40 [2464]);
assign l_39[1441]    = ( l_40 [2465]);
assign l_39[1442]    = ( l_40 [2466]);
assign l_39[1443]    = ( l_40 [2467]);
assign l_39[1444]    = ( l_40 [2468]);
assign l_39[1445]    = ( l_40 [2469]);
assign l_39[1446]    = ( l_40 [2470]);
assign l_39[1447]    = ( l_40 [2471]);
assign l_39[1448]    = ( l_40 [2472]);
assign l_39[1449]    = ( l_40 [2473]);
assign l_39[1450]    = ( l_40 [2474]);
assign l_39[1451]    = ( l_40 [2475]);
assign l_39[1452]    = ( l_40 [2476]);
assign l_39[1453]    = ( l_40 [2477]);
assign l_39[1454]    = ( l_40 [2478]);
assign l_39[1455]    = ( l_40 [2479]);
assign l_39[1456]    = ( l_40 [2480]);
assign l_39[1457]    = ( l_40 [2481]);
assign l_39[1458]    = ( l_40 [2482]);
assign l_39[1459]    = ( l_40 [2483]);
assign l_39[1460]    = ( l_40 [2484]);
assign l_39[1461]    = ( l_40 [2485]);
assign l_39[1462]    = ( l_40 [2486]);
assign l_39[1463]    = ( l_40 [2487]);
assign l_39[1464]    = ( l_40 [2488]);
assign l_39[1465]    = ( l_40 [2489]);
assign l_39[1466]    = ( l_40 [2490]);
assign l_39[1467]    = ( l_40 [2491]);
assign l_39[1468]    = ( l_40 [2492]);
assign l_39[1469]    = ( l_40 [2493]);
assign l_39[1470]    = ( l_40 [2494]);
assign l_39[1471]    = ( l_40 [2495]);
assign l_39[1472]    = ( l_40 [2496]);
assign l_39[1473]    = ( l_40 [2497]);
assign l_39[1474]    = ( l_40 [2498]);
assign l_39[1475]    = ( l_40 [2499]);
assign l_39[1476]    = ( l_40 [2500]);
assign l_39[1477]    = ( l_40 [2501]);
assign l_39[1478]    = ( l_40 [2502]);
assign l_39[1479]    = ( l_40 [2503]);
assign l_39[1480]    = ( l_40 [2504]);
assign l_39[1481]    = ( l_40 [2505]);
assign l_39[1482]    = ( l_40 [2506]);
assign l_39[1483]    = ( l_40 [2507]);
assign l_39[1484]    = ( l_40 [2508]);
assign l_39[1485]    = ( l_40 [2509]);
assign l_39[1486]    = ( l_40 [2510]);
assign l_39[1487]    = ( l_40 [2511]);
assign l_39[1488]    = ( l_40 [2512]);
assign l_39[1489]    = ( l_40 [2513]);
assign l_39[1490]    = ( l_40 [2514]);
assign l_39[1491]    = ( l_40 [2515]);
assign l_39[1492]    = ( l_40 [2516]);
assign l_39[1493]    = ( l_40 [2517]);
assign l_39[1494]    = ( l_40 [2518]);
assign l_39[1495]    = ( l_40 [2519]);
assign l_39[1496]    = ( l_40 [2520]);
assign l_39[1497]    = ( l_40 [2521]);
assign l_39[1498]    = ( l_40 [2522]);
assign l_39[1499]    = ( l_40 [2523]);
assign l_39[1500]    = ( l_40 [2524]);
assign l_39[1501]    = ( l_40 [2525]);
assign l_39[1502]    = ( l_40 [2526]);
assign l_39[1503]    = ( l_40 [2527]);
assign l_39[1504]    = ( l_40 [2528]);
assign l_39[1505]    = ( l_40 [2529]);
assign l_39[1506]    = ( l_40 [2530]);
assign l_39[1507]    = ( l_40 [2531]);
assign l_39[1508]    = ( l_40 [2532]);
assign l_39[1509]    = ( l_40 [2533]);
assign l_39[1510]    = ( l_40 [2534]);
assign l_39[1511]    = ( l_40 [2535]);
assign l_39[1512]    = ( l_40 [2536]);
assign l_39[1513]    = ( l_40 [2537]);
assign l_39[1514]    = ( l_40 [2538]);
assign l_39[1515]    = ( l_40 [2539]);
assign l_39[1516]    = ( l_40 [2540]);
assign l_39[1517]    = ( l_40 [2541]);
assign l_39[1518]    = ( l_40 [2542]);
assign l_39[1519]    = ( l_40 [2543]);
assign l_39[1520]    = ( l_40 [2544]);
assign l_39[1521]    = ( l_40 [2545]);
assign l_39[1522]    = ( l_40 [2546]);
assign l_39[1523]    = ( l_40 [2547]);
assign l_39[1524]    = ( l_40 [2548]);
assign l_39[1525]    = ( l_40 [2549]);
assign l_39[1526]    = ( l_40 [2550]);
assign l_39[1527]    = ( l_40 [2551]);
assign l_39[1528]    = ( l_40 [2552]);
assign l_39[1529]    = ( l_40 [2553]);
assign l_39[1530]    = ( l_40 [2554]);
assign l_39[1531]    = ( l_40 [2555]);
assign l_39[1532]    = ( l_40 [2556]);
assign l_39[1533]    = ( l_40 [2557]);
assign l_39[1534]    = ( l_40 [2558]);
assign l_39[1535]    = ( l_40 [2559]);
assign l_39[1536]    = ( l_40 [2560]);
assign l_39[1537]    = ( l_40 [2561]);
assign l_39[1538]    = ( l_40 [2562]);
assign l_39[1539]    = ( l_40 [2563]);
assign l_39[1540]    = ( l_40 [2564]);
assign l_39[1541]    = ( l_40 [2565]);
assign l_39[1542]    = ( l_40 [2566]);
assign l_39[1543]    = ( l_40 [2567]);
assign l_39[1544]    = ( l_40 [2568]);
assign l_39[1545]    = ( l_40 [2569]);
assign l_39[1546]    = ( l_40 [2570]);
assign l_39[1547]    = ( l_40 [2571]);
assign l_39[1548]    = ( l_40 [2572]);
assign l_39[1549]    = ( l_40 [2573]);
assign l_39[1550]    = ( l_40 [2574]);
assign l_39[1551]    = ( l_40 [2575]);
assign l_39[1552]    = ( l_40 [2576]);
assign l_39[1553]    = ( l_40 [2577]);
assign l_39[1554]    = ( l_40 [2578]);
assign l_39[1555]    = ( l_40 [2579]);
assign l_39[1556]    = ( l_40 [2580]);
assign l_39[1557]    = ( l_40 [2581]);
assign l_39[1558]    = ( l_40 [2582]);
assign l_39[1559]    = ( l_40 [2583]);
assign l_39[1560]    = ( l_40 [2584]);
assign l_39[1561]    = ( l_40 [2585]);
assign l_39[1562]    = ( l_40 [2586]);
assign l_39[1563]    = ( l_40 [2587]);
assign l_39[1564]    = ( l_40 [2588]);
assign l_39[1565]    = ( l_40 [2589]);
assign l_39[1566]    = ( l_40 [2590]);
assign l_39[1567]    = ( l_40 [2591]);
assign l_39[1568]    = ( l_40 [2592]);
assign l_39[1569]    = ( l_40 [2593]);
assign l_39[1570]    = ( l_40 [2594]);
assign l_39[1571]    = ( l_40 [2595]);
assign l_39[1572]    = ( l_40 [2596]);
assign l_39[1573]    = ( l_40 [2597]);
assign l_39[1574]    = ( l_40 [2598]);
assign l_39[1575]    = ( l_40 [2599]);
assign l_39[1576]    = ( l_40 [2600]);
assign l_39[1577]    = ( l_40 [2601]);
assign l_39[1578]    = ( l_40 [2602]);
assign l_39[1579]    = ( l_40 [2603]);
assign l_39[1580]    = ( l_40 [2604]);
assign l_39[1581]    = ( l_40 [2605]);
assign l_39[1582]    = ( l_40 [2606]);
assign l_39[1583]    = ( l_40 [2607]);
assign l_39[1584]    = ( l_40 [2608]);
assign l_39[1585]    = ( l_40 [2609]);
assign l_39[1586]    = ( l_40 [2610]);
assign l_39[1587]    = ( l_40 [2611]);
assign l_39[1588]    = ( l_40 [2612]);
assign l_39[1589]    = ( l_40 [2613]);
assign l_39[1590]    = ( l_40 [2614]);
assign l_39[1591]    = ( l_40 [2615]);
assign l_39[1592]    = ( l_40 [2616]);
assign l_39[1593]    = ( l_40 [2617]);
assign l_39[1594]    = ( l_40 [2618]);
assign l_39[1595]    = ( l_40 [2619]);
assign l_39[1596]    = ( l_40 [2620]);
assign l_39[1597]    = ( l_40 [2621]);
assign l_39[1598]    = ( l_40 [2622]);
assign l_39[1599]    = ( l_40 [2623]);
assign l_39[1600]    = ( l_40 [2624]);
assign l_39[1601]    = ( l_40 [2625]);
assign l_39[1602]    = ( l_40 [2626]);
assign l_39[1603]    = ( l_40 [2627]);
assign l_39[1604]    = ( l_40 [2628]);
assign l_39[1605]    = ( l_40 [2629]);
assign l_39[1606]    = ( l_40 [2630]);
assign l_39[1607]    = ( l_40 [2631]);
assign l_39[1608]    = ( l_40 [2632]);
assign l_39[1609]    = ( l_40 [2633]);
assign l_39[1610]    = ( l_40 [2634]);
assign l_39[1611]    = ( l_40 [2635]);
assign l_39[1612]    = ( l_40 [2636]);
assign l_39[1613]    = ( l_40 [2637]);
assign l_39[1614]    = ( l_40 [2638]);
assign l_39[1615]    = ( l_40 [2639]);
assign l_39[1616]    = ( l_40 [2640]);
assign l_39[1617]    = ( l_40 [2641]);
assign l_39[1618]    = ( l_40 [2642]);
assign l_39[1619]    = ( l_40 [2643]);
assign l_39[1620]    = ( l_40 [2644]);
assign l_39[1621]    = ( l_40 [2645]);
assign l_39[1622]    = ( l_40 [2646]);
assign l_39[1623]    = ( l_40 [2647]);
assign l_39[1624]    = ( l_40 [2648]);
assign l_39[1625]    = ( l_40 [2649]);
assign l_39[1626]    = ( l_40 [2650]);
assign l_39[1627]    = ( l_40 [2651]);
assign l_39[1628]    = ( l_40 [2652]);
assign l_39[1629]    = ( l_40 [2653]);
assign l_39[1630]    = ( l_40 [2654]);
assign l_39[1631]    = ( l_40 [2655]);
assign l_39[1632]    = ( l_40 [2656]);
assign l_39[1633]    = ( l_40 [2657]);
assign l_39[1634]    = ( l_40 [2658]);
assign l_39[1635]    = ( l_40 [2659]);
assign l_39[1636]    = ( l_40 [2660]);
assign l_39[1637]    = ( l_40 [2661]);
assign l_39[1638]    = ( l_40 [2662]);
assign l_39[1639]    = ( l_40 [2663]);
assign l_39[1640]    = ( l_40 [2664]);
assign l_39[1641]    = ( l_40 [2665]);
assign l_39[1642]    = ( l_40 [2666]);
assign l_39[1643]    = ( l_40 [2667]);
assign l_39[1644]    = ( l_40 [2668]);
assign l_39[1645]    = ( l_40 [2669]);
assign l_39[1646]    = ( l_40 [2670]);
assign l_39[1647]    = ( l_40 [2671]);
assign l_39[1648]    = ( l_40 [2672]);
assign l_39[1649]    = ( l_40 [2673]);
assign l_39[1650]    = ( l_40 [2674]);
assign l_39[1651]    = ( l_40 [2675]);
assign l_39[1652]    = ( l_40 [2676]);
assign l_39[1653]    = ( l_40 [2677]);
assign l_39[1654]    = ( l_40 [2678]);
assign l_39[1655]    = ( l_40 [2679]);
assign l_39[1656]    = ( l_40 [2680]);
assign l_39[1657]    = ( l_40 [2681]);
assign l_39[1658]    = ( l_40 [2682]);
assign l_39[1659]    = ( l_40 [2683]);
assign l_39[1660]    = ( l_40 [2684]);
assign l_39[1661]    = ( l_40 [2685]);
assign l_39[1662]    = ( l_40 [2686]);
assign l_39[1663]    = ( l_40 [2687]);
assign l_39[1664]    = ( l_40 [2688]);
assign l_39[1665]    = ( l_40 [2689]);
assign l_39[1666]    = ( l_40 [2690]);
assign l_39[1667]    = ( l_40 [2691]);
assign l_39[1668]    = ( l_40 [2692]);
assign l_39[1669]    = ( l_40 [2693]);
assign l_39[1670]    = ( l_40 [2694]);
assign l_39[1671]    = ( l_40 [2695]);
assign l_39[1672]    = ( l_40 [2696]);
assign l_39[1673]    = ( l_40 [2697]);
assign l_39[1674]    = ( l_40 [2698]);
assign l_39[1675]    = ( l_40 [2699]);
assign l_39[1676]    = ( l_40 [2700]);
assign l_39[1677]    = ( l_40 [2701]);
assign l_39[1678]    = ( l_40 [2702]);
assign l_39[1679]    = ( l_40 [2703]);
assign l_39[1680]    = ( l_40 [2704]);
assign l_39[1681]    = ( l_40 [2705]);
assign l_39[1682]    = ( l_40 [2706]);
assign l_39[1683]    = ( l_40 [2707]);
assign l_39[1684]    = ( l_40 [2708]);
assign l_39[1685]    = ( l_40 [2709]);
assign l_39[1686]    = ( l_40 [2710]);
assign l_39[1687]    = ( l_40 [2711]);
assign l_39[1688]    = ( l_40 [2712]);
assign l_39[1689]    = ( l_40 [2713]);
assign l_39[1690]    = ( l_40 [2714]);
assign l_39[1691]    = ( l_40 [2715]);
assign l_39[1692]    = ( l_40 [2716]);
assign l_39[1693]    = ( l_40 [2717]);
assign l_39[1694]    = ( l_40 [2718]);
assign l_39[1695]    = ( l_40 [2719]);
assign l_39[1696]    = ( l_40 [2720]);
assign l_39[1697]    = ( l_40 [2721]);
assign l_39[1698]    = ( l_40 [2722]);
assign l_39[1699]    = ( l_40 [2723]);
assign l_39[1700]    = ( l_40 [2724]);
assign l_39[1701]    = ( l_40 [2725]);
assign l_39[1702]    = ( l_40 [2726]);
assign l_39[1703]    = ( l_40 [2727]);
assign l_39[1704]    = ( l_40 [2728]);
assign l_39[1705]    = ( l_40 [2729]);
assign l_39[1706]    = ( l_40 [2730]);
assign l_39[1707]    = ( l_40 [2731]);
assign l_39[1708]    = ( l_40 [2732]);
assign l_39[1709]    = ( l_40 [2733]);
assign l_39[1710]    = ( l_40 [2734]);
assign l_39[1711]    = ( l_40 [2735]);
assign l_39[1712]    = ( l_40 [2736]);
assign l_39[1713]    = ( l_40 [2737]);
assign l_39[1714]    = ( l_40 [2738]);
assign l_39[1715]    = ( l_40 [2739]);
assign l_39[1716]    = ( l_40 [2740]);
assign l_39[1717]    = ( l_40 [2741]);
assign l_39[1718]    = ( l_40 [2742]);
assign l_39[1719]    = ( l_40 [2743]);
assign l_39[1720]    = ( l_40 [2744]);
assign l_39[1721]    = ( l_40 [2745]);
assign l_39[1722]    = ( l_40 [2746]);
assign l_39[1723]    = ( l_40 [2747]);
assign l_39[1724]    = ( l_40 [2748]);
assign l_39[1725]    = ( l_40 [2749]);
assign l_39[1726]    = ( l_40 [2750]);
assign l_39[1727]    = ( l_40 [2751]);
assign l_39[1728]    = ( l_40 [2752]);
assign l_39[1729]    = ( l_40 [2753]);
assign l_39[1730]    = ( l_40 [2754]);
assign l_39[1731]    = ( l_40 [2755]);
assign l_39[1732]    = ( l_40 [2756]);
assign l_39[1733]    = ( l_40 [2757]);
assign l_39[1734]    = ( l_40 [2758]);
assign l_39[1735]    = ( l_40 [2759]);
assign l_39[1736]    = ( l_40 [2760]);
assign l_39[1737]    = ( l_40 [2761]);
assign l_39[1738]    = ( l_40 [2762]);
assign l_39[1739]    = ( l_40 [2763]);
assign l_39[1740]    = ( l_40 [2764]);
assign l_39[1741]    = ( l_40 [2765]);
assign l_39[1742]    = ( l_40 [2766]);
assign l_39[1743]    = ( l_40 [2767]);
assign l_39[1744]    = ( l_40 [2768]);
assign l_39[1745]    = ( l_40 [2769]);
assign l_39[1746]    = ( l_40 [2770]);
assign l_39[1747]    = ( l_40 [2771]);
assign l_39[1748]    = ( l_40 [2772]);
assign l_39[1749]    = ( l_40 [2773]);
assign l_39[1750]    = ( l_40 [2774]);
assign l_39[1751]    = ( l_40 [2775]);
assign l_39[1752]    = ( l_40 [2776]);
assign l_39[1753]    = ( l_40 [2777]);
assign l_39[1754]    = ( l_40 [2778]);
assign l_39[1755]    = ( l_40 [2779]);
assign l_39[1756]    = ( l_40 [2780]);
assign l_39[1757]    = ( l_40 [2781]);
assign l_39[1758]    = ( l_40 [2782]);
assign l_39[1759]    = ( l_40 [2783]);
assign l_39[1760]    = ( l_40 [2784]);
assign l_39[1761]    = ( l_40 [2785]);
assign l_39[1762]    = ( l_40 [2786]);
assign l_39[1763]    = ( l_40 [2787]);
assign l_39[1764]    = ( l_40 [2788]);
assign l_39[1765]    = ( l_40 [2789]);
assign l_39[1766]    = ( l_40 [2790]);
assign l_39[1767]    = ( l_40 [2791]);
assign l_39[1768]    = ( l_40 [2792]);
assign l_39[1769]    = ( l_40 [2793]);
assign l_39[1770]    = ( l_40 [2794]);
assign l_39[1771]    = ( l_40 [2795]);
assign l_39[1772]    = ( l_40 [2796]);
assign l_39[1773]    = ( l_40 [2797]);
assign l_39[1774]    = ( l_40 [2798]);
assign l_39[1775]    = ( l_40 [2799]);
assign l_39[1776]    = ( l_40 [2800]);
assign l_39[1777]    = ( l_40 [2801]);
assign l_39[1778]    = ( l_40 [2802]);
assign l_39[1779]    = ( l_40 [2803]);
assign l_39[1780]    = ( l_40 [2804]);
assign l_39[1781]    = ( l_40 [2805]);
assign l_39[1782]    = ( l_40 [2806]);
assign l_39[1783]    = ( l_40 [2807]);
assign l_39[1784]    = ( l_40 [2808]);
assign l_39[1785]    = ( l_40 [2809]);
assign l_39[1786]    = ( l_40 [2810]);
assign l_39[1787]    = ( l_40 [2811]);
assign l_39[1788]    = ( l_40 [2812]);
assign l_39[1789]    = ( l_40 [2813]);
assign l_39[1790]    = ( l_40 [2814]);
assign l_39[1791]    = ( l_40 [2815]);
assign l_39[1792]    = ( l_40 [2816]);
assign l_39[1793]    = ( l_40 [2817]);
assign l_39[1794]    = ( l_40 [2818]);
assign l_39[1795]    = ( l_40 [2819]);
assign l_39[1796]    = ( l_40 [2820]);
assign l_39[1797]    = ( l_40 [2821]);
assign l_39[1798]    = ( l_40 [2822]);
assign l_39[1799]    = ( l_40 [2823]);
assign l_39[1800]    = ( l_40 [2824]);
assign l_39[1801]    = ( l_40 [2825]);
assign l_39[1802]    = ( l_40 [2826]);
assign l_39[1803]    = ( l_40 [2827]);
assign l_39[1804]    = ( l_40 [2828]);
assign l_39[1805]    = ( l_40 [2829]);
assign l_39[1806]    = ( l_40 [2830]);
assign l_39[1807]    = ( l_40 [2831]);
assign l_39[1808]    = ( l_40 [2832]);
assign l_39[1809]    = ( l_40 [2833]);
assign l_39[1810]    = ( l_40 [2834]);
assign l_39[1811]    = ( l_40 [2835]);
assign l_39[1812]    = ( l_40 [2836]);
assign l_39[1813]    = ( l_40 [2837]);
assign l_39[1814]    = ( l_40 [2838]);
assign l_39[1815]    = ( l_40 [2839]);
assign l_39[1816]    = ( l_40 [2840]);
assign l_39[1817]    = ( l_40 [2841]);
assign l_39[1818]    = ( l_40 [2842]);
assign l_39[1819]    = ( l_40 [2843]);
assign l_39[1820]    = ( l_40 [2844]);
assign l_39[1821]    = ( l_40 [2845]);
assign l_39[1822]    = ( l_40 [2846]);
assign l_39[1823]    = ( l_40 [2847]);
assign l_39[1824]    = ( l_40 [2848]);
assign l_39[1825]    = ( l_40 [2849]);
assign l_39[1826]    = ( l_40 [2850]);
assign l_39[1827]    = ( l_40 [2851]);
assign l_39[1828]    = ( l_40 [2852]);
assign l_39[1829]    = ( l_40 [2853]);
assign l_39[1830]    = ( l_40 [2854]);
assign l_39[1831]    = ( l_40 [2855]);
assign l_39[1832]    = ( l_40 [2856]);
assign l_39[1833]    = ( l_40 [2857]);
assign l_39[1834]    = ( l_40 [2858]);
assign l_39[1835]    = ( l_40 [2859]);
assign l_39[1836]    = ( l_40 [2860]);
assign l_39[1837]    = ( l_40 [2861]);
assign l_39[1838]    = ( l_40 [2862]);
assign l_39[1839]    = ( l_40 [2863]);
assign l_39[1840]    = ( l_40 [2864]);
assign l_39[1841]    = ( l_40 [2865]);
assign l_39[1842]    = ( l_40 [2866]);
assign l_39[1843]    = ( l_40 [2867]);
assign l_39[1844]    = ( l_40 [2868]);
assign l_39[1845]    = ( l_40 [2869]);
assign l_39[1846]    = ( l_40 [2870]);
assign l_39[1847]    = ( l_40 [2871]);
assign l_39[1848]    = ( l_40 [2872]);
assign l_39[1849]    = ( l_40 [2873]);
assign l_39[1850]    = ( l_40 [2874]);
assign l_39[1851]    = ( l_40 [2875]);
assign l_39[1852]    = ( l_40 [2876]);
assign l_39[1853]    = ( l_40 [2877]);
assign l_39[1854]    = ( l_40 [2878]);
assign l_39[1855]    = ( l_40 [2879]);
assign l_39[1856]    = ( l_40 [2880]);
assign l_39[1857]    = ( l_40 [2881]);
assign l_39[1858]    = ( l_40 [2882]);
assign l_39[1859]    = ( l_40 [2883]);
assign l_39[1860]    = ( l_40 [2884]);
assign l_39[1861]    = ( l_40 [2885]);
assign l_39[1862]    = ( l_40 [2886]);
assign l_39[1863]    = ( l_40 [2887]);
assign l_39[1864]    = ( l_40 [2888]);
assign l_39[1865]    = ( l_40 [2889]);
assign l_39[1866]    = ( l_40 [2890]);
assign l_39[1867]    = ( l_40 [2891]);
assign l_39[1868]    = ( l_40 [2892]);
assign l_39[1869]    = ( l_40 [2893]);
assign l_39[1870]    = ( l_40 [2894]);
assign l_39[1871]    = ( l_40 [2895]);
assign l_39[1872]    = ( l_40 [2896]);
assign l_39[1873]    = ( l_40 [2897]);
assign l_39[1874]    = ( l_40 [2898]);
assign l_39[1875]    = ( l_40 [2899]);
assign l_39[1876]    = ( l_40 [2900]);
assign l_39[1877]    = ( l_40 [2901]);
assign l_39[1878]    = ( l_40 [2902]);
assign l_39[1879]    = ( l_40 [2903]);
assign l_39[1880]    = ( l_40 [2904]);
assign l_39[1881]    = ( l_40 [2905]);
assign l_39[1882]    = ( l_40 [2906]);
assign l_39[1883]    = ( l_40 [2907]);
assign l_39[1884]    = ( l_40 [2908]);
assign l_39[1885]    = ( l_40 [2909]);
assign l_39[1886]    = ( l_40 [2910]);
assign l_39[1887]    = ( l_40 [2911]);
assign l_39[1888]    = ( l_40 [2912]);
assign l_39[1889]    = ( l_40 [2913]);
assign l_39[1890]    = ( l_40 [2914]);
assign l_39[1891]    = ( l_40 [2915]);
assign l_39[1892]    = ( l_40 [2916]);
assign l_39[1893]    = ( l_40 [2917]);
assign l_39[1894]    = ( l_40 [2918]);
assign l_39[1895]    = ( l_40 [2919]);
assign l_39[1896]    = ( l_40 [2920]);
assign l_39[1897]    = ( l_40 [2921]);
assign l_39[1898]    = ( l_40 [2922]);
assign l_39[1899]    = ( l_40 [2923]);
assign l_39[1900]    = ( l_40 [2924]);
assign l_39[1901]    = ( l_40 [2925]);
assign l_39[1902]    = ( l_40 [2926]);
assign l_39[1903]    = ( l_40 [2927]);
assign l_39[1904]    = ( l_40 [2928]);
assign l_39[1905]    = ( l_40 [2929]);
assign l_39[1906]    = ( l_40 [2930]);
assign l_39[1907]    = ( l_40 [2931]);
assign l_39[1908]    = ( l_40 [2932]);
assign l_39[1909]    = ( l_40 [2933]);
assign l_39[1910]    = ( l_40 [2934]);
assign l_39[1911]    = ( l_40 [2935]);
assign l_39[1912]    = ( l_40 [2936]);
assign l_39[1913]    = ( l_40 [2937]);
assign l_39[1914]    = ( l_40 [2938]);
assign l_39[1915]    = ( l_40 [2939]);
assign l_39[1916]    = ( l_40 [2940]);
assign l_39[1917]    = ( l_40 [2941]);
assign l_39[1918]    = ( l_40 [2942]);
assign l_39[1919]    = ( l_40 [2943]);
assign l_39[1920]    = ( l_40 [2944]);
assign l_39[1921]    = ( l_40 [2945]);
assign l_39[1922]    = ( l_40 [2946]);
assign l_39[1923]    = ( l_40 [2947]);
assign l_39[1924]    = ( l_40 [2948]);
assign l_39[1925]    = ( l_40 [2949]);
assign l_39[1926]    = ( l_40 [2950]);
assign l_39[1927]    = ( l_40 [2951]);
assign l_39[1928]    = ( l_40 [2952]);
assign l_39[1929]    = ( l_40 [2953]);
assign l_39[1930]    = ( l_40 [2954]);
assign l_39[1931]    = ( l_40 [2955]);
assign l_39[1932]    = ( l_40 [2956]);
assign l_39[1933]    = ( l_40 [2957]);
assign l_39[1934]    = ( l_40 [2958]);
assign l_39[1935]    = ( l_40 [2959]);
assign l_39[1936]    = ( l_40 [2960]);
assign l_39[1937]    = ( l_40 [2961]);
assign l_39[1938]    = ( l_40 [2962]);
assign l_39[1939]    = ( l_40 [2963]);
assign l_39[1940]    = ( l_40 [2964]);
assign l_39[1941]    = ( l_40 [2965]);
assign l_39[1942]    = ( l_40 [2966]);
assign l_39[1943]    = ( l_40 [2967]);
assign l_39[1944]    = ( l_40 [2968]);
assign l_39[1945]    = ( l_40 [2969]);
assign l_39[1946]    = ( l_40 [2970]);
assign l_39[1947]    = ( l_40 [2971]);
assign l_39[1948]    = ( l_40 [2972]);
assign l_39[1949]    = ( l_40 [2973]);
assign l_39[1950]    = ( l_40 [2974]);
assign l_39[1951]    = ( l_40 [2975]);
assign l_39[1952]    = ( l_40 [2976]);
assign l_39[1953]    = ( l_40 [2977]);
assign l_39[1954]    = ( l_40 [2978]);
assign l_39[1955]    = ( l_40 [2979]);
assign l_39[1956]    = ( l_40 [2980]);
assign l_39[1957]    = ( l_40 [2981]);
assign l_39[1958]    = ( l_40 [2982]);
assign l_39[1959]    = ( l_40 [2983]);
assign l_39[1960]    = ( l_40 [2984]);
assign l_39[1961]    = ( l_40 [2985]);
assign l_39[1962]    = ( l_40 [2986]);
assign l_39[1963]    = ( l_40 [2987]);
assign l_39[1964]    = ( l_40 [2988]);
assign l_39[1965]    = ( l_40 [2989]);
assign l_39[1966]    = ( l_40 [2990]);
assign l_39[1967]    = ( l_40 [2991]);
assign l_39[1968]    = ( l_40 [2992]);
assign l_39[1969]    = ( l_40 [2993]);
assign l_39[1970]    = ( l_40 [2994]);
assign l_39[1971]    = ( l_40 [2995]);
assign l_39[1972]    = ( l_40 [2996]);
assign l_39[1973]    = ( l_40 [2997]);
assign l_39[1974]    = ( l_40 [2998]);
assign l_39[1975]    = ( l_40 [2999]);
assign l_39[1976]    = ( l_40 [3000]);
assign l_39[1977]    = ( l_40 [3001]);
assign l_39[1978]    = ( l_40 [3002]);
assign l_39[1979]    = ( l_40 [3003]);
assign l_39[1980]    = ( l_40 [3004]);
assign l_39[1981]    = ( l_40 [3005]);
assign l_39[1982]    = ( l_40 [3006]);
assign l_39[1983]    = ( l_40 [3007]);
assign l_39[1984]    = ( l_40 [3008]);
assign l_39[1985]    = ( l_40 [3009]);
assign l_39[1986]    = ( l_40 [3010]);
assign l_39[1987]    = ( l_40 [3011]);
assign l_39[1988]    = ( l_40 [3012]);
assign l_39[1989]    = ( l_40 [3013]);
assign l_39[1990]    = ( l_40 [3014]);
assign l_39[1991]    = ( l_40 [3015]);
assign l_39[1992]    = ( l_40 [3016]);
assign l_39[1993]    = ( l_40 [3017]);
assign l_39[1994]    = ( l_40 [3018]);
assign l_39[1995]    = ( l_40 [3019]);
assign l_39[1996]    = ( l_40 [3020]);
assign l_39[1997]    = ( l_40 [3021]);
assign l_39[1998]    = ( l_40 [3022]);
assign l_39[1999]    = ( l_40 [3023]);
assign l_39[2000]    = ( l_40 [3024]);
assign l_39[2001]    = ( l_40 [3025]);
assign l_39[2002]    = ( l_40 [3026]);
assign l_39[2003]    = ( l_40 [3027]);
assign l_39[2004]    = ( l_40 [3028]);
assign l_39[2005]    = ( l_40 [3029]);
assign l_39[2006]    = ( l_40 [3030]);
assign l_39[2007]    = ( l_40 [3031]);
assign l_39[2008]    = ( l_40 [3032]);
assign l_39[2009]    = ( l_40 [3033]);
assign l_39[2010]    = ( l_40 [3034]);
assign l_39[2011]    = ( l_40 [3035]);
assign l_39[2012]    = ( l_40 [3036]);
assign l_39[2013]    = ( l_40 [3037]);
assign l_39[2014]    = ( l_40 [3038]);
assign l_39[2015]    = ( l_40 [3039]);
assign l_39[2016]    = ( l_40 [3040]);
assign l_39[2017]    = ( l_40 [3041]);
assign l_39[2018]    = ( l_40 [3042]);
assign l_39[2019]    = ( l_40 [3043]);
assign l_39[2020]    = ( l_40 [3044]);
assign l_39[2021]    = ( l_40 [3045]);
assign l_39[2022]    = ( l_40 [3046]);
assign l_39[2023]    = ( l_40 [3047]);
assign l_39[2024]    = ( l_40 [3048]);
assign l_39[2025]    = ( l_40 [3049]);
assign l_39[2026]    = ( l_40 [3050]);
assign l_39[2027]    = ( l_40 [3051]);
assign l_39[2028]    = ( l_40 [3052]);
assign l_39[2029]    = ( l_40 [3053]);
assign l_39[2030]    = ( l_40 [3054]);
assign l_39[2031]    = ( l_40 [3055]);
assign l_39[2032]    = ( l_40 [3056]);
assign l_39[2033]    = ( l_40 [3057]);
assign l_39[2034]    = ( l_40 [3058]);
assign l_39[2035]    = ( l_40 [3059]);
assign l_39[2036]    = ( l_40 [3060]);
assign l_39[2037]    = ( l_40 [3061]);
assign l_39[2038]    = ( l_40 [3062]);
assign l_39[2039]    = ( l_40 [3063]);
assign l_39[2040]    = ( l_40 [3064]);
assign l_39[2041]    = ( l_40 [3065]);
assign l_39[2042]    = ( l_40 [3066]);
assign l_39[2043]    = ( l_40 [3067]);
assign l_39[2044]    = ( l_40 [3068]);
assign l_39[2045]    = ( l_40 [3069]);
assign l_39[2046]    = ( l_40 [3070]);
assign l_39[2047]    = ( l_40 [3071]);
assign l_39[2048]    = ( l_40 [3072]);
assign l_39[2049]    = ( l_40 [3073]);
assign l_39[2050]    = ( l_40 [3074]);
assign l_39[2051]    = ( l_40 [3075]);
assign l_39[2052]    = ( l_40 [3076]);
assign l_39[2053]    = ( l_40 [3077]);
assign l_39[2054]    = ( l_40 [3078]);
assign l_39[2055]    = ( l_40 [3079]);
assign l_39[2056]    = ( l_40 [3080]);
assign l_39[2057]    = ( l_40 [3081]);
assign l_39[2058]    = ( l_40 [3082]);
assign l_39[2059]    = ( l_40 [3083]);
assign l_39[2060]    = ( l_40 [3084]);
assign l_39[2061]    = ( l_40 [3085]);
assign l_39[2062]    = ( l_40 [3086]);
assign l_39[2063]    = ( l_40 [3087]);
assign l_39[2064]    = ( l_40 [3088]);
assign l_39[2065]    = ( l_40 [3089]);
assign l_39[2066]    = ( l_40 [3090]);
assign l_39[2067]    = ( l_40 [3091]);
assign l_39[2068]    = ( l_40 [3092]);
assign l_39[2069]    = ( l_40 [3093]);
assign l_39[2070]    = ( l_40 [3094]);
assign l_39[2071]    = ( l_40 [3095]);
assign l_39[2072]    = ( l_40 [3096]);
assign l_39[2073]    = ( l_40 [3097]);
assign l_39[2074]    = ( l_40 [3098]);
assign l_39[2075]    = ( l_40 [3099]);
assign l_39[2076]    = ( l_40 [3100]);
assign l_39[2077]    = ( l_40 [3101]);
assign l_39[2078]    = ( l_40 [3102]);
assign l_39[2079]    = ( l_40 [3103]);
assign l_39[2080]    = ( l_40 [3104]);
assign l_39[2081]    = ( l_40 [3105]);
assign l_39[2082]    = ( l_40 [3106]);
assign l_39[2083]    = ( l_40 [3107]);
assign l_39[2084]    = ( l_40 [3108]);
assign l_39[2085]    = ( l_40 [3109]);
assign l_39[2086]    = ( l_40 [3110]);
assign l_39[2087]    = ( l_40 [3111]);
assign l_39[2088]    = ( l_40 [3112]);
assign l_39[2089]    = ( l_40 [3113]);
assign l_39[2090]    = ( l_40 [3114]);
assign l_39[2091]    = ( l_40 [3115]);
assign l_39[2092]    = ( l_40 [3116]);
assign l_39[2093]    = ( l_40 [3117]);
assign l_39[2094]    = ( l_40 [3118]);
assign l_39[2095]    = ( l_40 [3119]);
assign l_39[2096]    = ( l_40 [3120]);
assign l_39[2097]    = ( l_40 [3121]);
assign l_39[2098]    = ( l_40 [3122]);
assign l_39[2099]    = ( l_40 [3123]);
assign l_39[2100]    = ( l_40 [3124]);
assign l_39[2101]    = ( l_40 [3125]);
assign l_39[2102]    = ( l_40 [3126]);
assign l_39[2103]    = ( l_40 [3127]);
assign l_39[2104]    = ( l_40 [3128]);
assign l_39[2105]    = ( l_40 [3129]);
assign l_39[2106]    = ( l_40 [3130]);
assign l_39[2107]    = ( l_40 [3131]);
assign l_39[2108]    = ( l_40 [3132]);
assign l_39[2109]    = ( l_40 [3133]);
assign l_39[2110]    = ( l_40 [3134]);
assign l_39[2111]    = ( l_40 [3135]);
assign l_39[2112]    = ( l_40 [3136]);
assign l_39[2113]    = ( l_40 [3137]);
assign l_39[2114]    = ( l_40 [3138]);
assign l_39[2115]    = ( l_40 [3139]);
assign l_39[2116]    = ( l_40 [3140]);
assign l_39[2117]    = ( l_40 [3141]);
assign l_39[2118]    = ( l_40 [3142]);
assign l_39[2119]    = ( l_40 [3143]);
assign l_39[2120]    = ( l_40 [3144]);
assign l_39[2121]    = ( l_40 [3145]);
assign l_39[2122]    = ( l_40 [3146]);
assign l_39[2123]    = ( l_40 [3147]);
assign l_39[2124]    = ( l_40 [3148]);
assign l_39[2125]    = ( l_40 [3149]);
assign l_39[2126]    = ( l_40 [3150]);
assign l_39[2127]    = ( l_40 [3151]);
assign l_39[2128]    = ( l_40 [3152]);
assign l_39[2129]    = ( l_40 [3153]);
assign l_39[2130]    = ( l_40 [3154]);
assign l_39[2131]    = ( l_40 [3155]);
assign l_39[2132]    = ( l_40 [3156]);
assign l_39[2133]    = ( l_40 [3157]);
assign l_39[2134]    = ( l_40 [3158]);
assign l_39[2135]    = ( l_40 [3159]);
assign l_39[2136]    = ( l_40 [3160]);
assign l_39[2137]    = ( l_40 [3161]);
assign l_39[2138]    = ( l_40 [3162]);
assign l_39[2139]    = ( l_40 [3163]);
assign l_39[2140]    = ( l_40 [3164]);
assign l_39[2141]    = ( l_40 [3165]);
assign l_39[2142]    = ( l_40 [3166]);
assign l_39[2143]    = ( l_40 [3167]);
assign l_39[2144]    = ( l_40 [3168]);
assign l_39[2145]    = ( l_40 [3169]);
assign l_39[2146]    = ( l_40 [3170]);
assign l_39[2147]    = ( l_40 [3171]);
assign l_39[2148]    = ( l_40 [3172]);
assign l_39[2149]    = ( l_40 [3173]);
assign l_39[2150]    = ( l_40 [3174]);
assign l_39[2151]    = ( l_40 [3175]);
assign l_39[2152]    = ( l_40 [3176]);
assign l_39[2153]    = ( l_40 [3177]);
assign l_39[2154]    = ( l_40 [3178]);
assign l_39[2155]    = ( l_40 [3179]);
assign l_39[2156]    = ( l_40 [3180]);
assign l_39[2157]    = ( l_40 [3181]);
assign l_39[2158]    = ( l_40 [3182]);
assign l_39[2159]    = ( l_40 [3183]);
assign l_39[2160]    = ( l_40 [3184]);
assign l_39[2161]    = ( l_40 [3185]);
assign l_39[2162]    = ( l_40 [3186]);
assign l_39[2163]    = ( l_40 [3187]);
assign l_39[2164]    = ( l_40 [3188]);
assign l_39[2165]    = ( l_40 [3189]);
assign l_39[2166]    = ( l_40 [3190]);
assign l_39[2167]    = ( l_40 [3191]);
assign l_39[2168]    = ( l_40 [3192]);
assign l_39[2169]    = ( l_40 [3193]);
assign l_39[2170]    = ( l_40 [3194]);
assign l_39[2171]    = ( l_40 [3195]);
assign l_39[2172]    = ( l_40 [3196]);
assign l_39[2173]    = ( l_40 [3197]);
assign l_39[2174]    = ( l_40 [3198]);
assign l_39[2175]    = ( l_40 [3199]);
assign l_39[2176]    = ( l_40 [3200]);
assign l_39[2177]    = ( l_40 [3201]);
assign l_39[2178]    = ( l_40 [3202]);
assign l_39[2179]    = ( l_40 [3203]);
assign l_39[2180]    = ( l_40 [3204]);
assign l_39[2181]    = ( l_40 [3205]);
assign l_39[2182]    = ( l_40 [3206]);
assign l_39[2183]    = ( l_40 [3207]);
assign l_39[2184]    = ( l_40 [3208]);
assign l_39[2185]    = ( l_40 [3209]);
assign l_39[2186]    = ( l_40 [3210]);
assign l_39[2187]    = ( l_40 [3211]);
assign l_39[2188]    = ( l_40 [3212]);
assign l_39[2189]    = ( l_40 [3213]);
assign l_39[2190]    = ( l_40 [3214]);
assign l_39[2191]    = ( l_40 [3215]);
assign l_39[2192]    = ( l_40 [3216]);
assign l_39[2193]    = ( l_40 [3217]);
assign l_39[2194]    = ( l_40 [3218]);
assign l_39[2195]    = ( l_40 [3219]);
assign l_39[2196]    = ( l_40 [3220]);
assign l_39[2197]    = ( l_40 [3221]);
assign l_39[2198]    = ( l_40 [3222]);
assign l_39[2199]    = ( l_40 [3223]);
assign l_39[2200]    = ( l_40 [3224]);
assign l_39[2201]    = ( l_40 [3225]);
assign l_39[2202]    = ( l_40 [3226]);
assign l_39[2203]    = ( l_40 [3227]);
assign l_39[2204]    = ( l_40 [3228]);
assign l_39[2205]    = ( l_40 [3229]);
assign l_39[2206]    = ( l_40 [3230]);
assign l_39[2207]    = ( l_40 [3231]);
assign l_39[2208]    = ( l_40 [3232]);
assign l_39[2209]    = ( l_40 [3233]);
assign l_39[2210]    = ( l_40 [3234]);
assign l_39[2211]    = ( l_40 [3235]);
assign l_39[2212]    = ( l_40 [3236]);
assign l_39[2213]    = ( l_40 [3237]);
assign l_39[2214]    = ( l_40 [3238]);
assign l_39[2215]    = ( l_40 [3239]);
assign l_39[2216]    = ( l_40 [3240]);
assign l_39[2217]    = ( l_40 [3241]);
assign l_39[2218]    = ( l_40 [3242]);
assign l_39[2219]    = ( l_40 [3243]);
assign l_39[2220]    = ( l_40 [3244]);
assign l_39[2221]    = ( l_40 [3245]);
assign l_39[2222]    = ( l_40 [3246]);
assign l_39[2223]    = ( l_40 [3247]);
assign l_39[2224]    = ( l_40 [3248]);
assign l_39[2225]    = ( l_40 [3249]);
assign l_39[2226]    = ( l_40 [3250]);
assign l_39[2227]    = ( l_40 [3251]);
assign l_39[2228]    = ( l_40 [3252]);
assign l_39[2229]    = ( l_40 [3253]);
assign l_39[2230]    = ( l_40 [3254]);
assign l_39[2231]    = ( l_40 [3255]);
assign l_39[2232]    = ( l_40 [3256]);
assign l_39[2233]    = ( l_40 [3257]);
assign l_39[2234]    = ( l_40 [3258]);
assign l_39[2235]    = ( l_40 [3259]);
assign l_39[2236]    = ( l_40 [3260]);
assign l_39[2237]    = ( l_40 [3261]);
assign l_39[2238]    = ( l_40 [3262]);
assign l_39[2239]    = ( l_40 [3263]);
assign l_39[2240]    = ( l_40 [3264]);
assign l_39[2241]    = ( l_40 [3265]);
assign l_39[2242]    = ( l_40 [3266]);
assign l_39[2243]    = ( l_40 [3267]);
assign l_39[2244]    = ( l_40 [3268]);
assign l_39[2245]    = ( l_40 [3269]);
assign l_39[2246]    = ( l_40 [3270]);
assign l_39[2247]    = ( l_40 [3271]);
assign l_39[2248]    = ( l_40 [3272]);
assign l_39[2249]    = ( l_40 [3273]);
assign l_39[2250]    = ( l_40 [3274]);
assign l_39[2251]    = ( l_40 [3275]);
assign l_39[2252]    = ( l_40 [3276]);
assign l_39[2253]    = ( l_40 [3277]);
assign l_39[2254]    = ( l_40 [3278]);
assign l_39[2255]    = ( l_40 [3279]);
assign l_39[2256]    = ( l_40 [3280]);
assign l_39[2257]    = ( l_40 [3281]);
assign l_39[2258]    = ( l_40 [3282]);
assign l_39[2259]    = ( l_40 [3283]);
assign l_39[2260]    = ( l_40 [3284]);
assign l_39[2261]    = ( l_40 [3285]);
assign l_39[2262]    = ( l_40 [3286]);
assign l_39[2263]    = ( l_40 [3287]);
assign l_39[2264]    = ( l_40 [3288]);
assign l_39[2265]    = ( l_40 [3289]);
assign l_39[2266]    = ( l_40 [3290]);
assign l_39[2267]    = ( l_40 [3291]);
assign l_39[2268]    = ( l_40 [3292]);
assign l_39[2269]    = ( l_40 [3293]);
assign l_39[2270]    = ( l_40 [3294]);
assign l_39[2271]    = ( l_40 [3295]);
assign l_39[2272]    = ( l_40 [3296]);
assign l_39[2273]    = ( l_40 [3297]);
assign l_39[2274]    = ( l_40 [3298]);
assign l_39[2275]    = ( l_40 [3299]);
assign l_39[2276]    = ( l_40 [3300]);
assign l_39[2277]    = ( l_40 [3301]);
assign l_39[2278]    = ( l_40 [3302]);
assign l_39[2279]    = ( l_40 [3303]);
assign l_39[2280]    = ( l_40 [3304]);
assign l_39[2281]    = ( l_40 [3305]);
assign l_39[2282]    = ( l_40 [3306]);
assign l_39[2283]    = ( l_40 [3307]);
assign l_39[2284]    = ( l_40 [3308]);
assign l_39[2285]    = ( l_40 [3309]);
assign l_39[2286]    = ( l_40 [3310]);
assign l_39[2287]    = ( l_40 [3311]);
assign l_39[2288]    = ( l_40 [3312]);
assign l_39[2289]    = ( l_40 [3313]);
assign l_39[2290]    = ( l_40 [3314]);
assign l_39[2291]    = ( l_40 [3315]);
assign l_39[2292]    = ( l_40 [3316]);
assign l_39[2293]    = ( l_40 [3317]);
assign l_39[2294]    = ( l_40 [3318]);
assign l_39[2295]    = ( l_40 [3319]);
assign l_39[2296]    = ( l_40 [3320]);
assign l_39[2297]    = ( l_40 [3321]);
assign l_39[2298]    = ( l_40 [3322]);
assign l_39[2299]    = ( l_40 [3323]);
assign l_39[2300]    = ( l_40 [3324]);
assign l_39[2301]    = ( l_40 [3325]);
assign l_39[2302]    = ( l_40 [3326]);
assign l_39[2303]    = ( l_40 [3327]);
assign l_39[2304]    = ( l_40 [3328]);
assign l_39[2305]    = ( l_40 [3329]);
assign l_39[2306]    = ( l_40 [3330]);
assign l_39[2307]    = ( l_40 [3331]);
assign l_39[2308]    = ( l_40 [3332]);
assign l_39[2309]    = ( l_40 [3333]);
assign l_39[2310]    = ( l_40 [3334]);
assign l_39[2311]    = ( l_40 [3335]);
assign l_39[2312]    = ( l_40 [3336]);
assign l_39[2313]    = ( l_40 [3337]);
assign l_39[2314]    = ( l_40 [3338]);
assign l_39[2315]    = ( l_40 [3339]);
assign l_39[2316]    = ( l_40 [3340]);
assign l_39[2317]    = ( l_40 [3341]);
assign l_39[2318]    = ( l_40 [3342]);
assign l_39[2319]    = ( l_40 [3343]);
assign l_39[2320]    = ( l_40 [3344]);
assign l_39[2321]    = ( l_40 [3345]);
assign l_39[2322]    = ( l_40 [3346]);
assign l_39[2323]    = ( l_40 [3347]);
assign l_39[2324]    = ( l_40 [3348]);
assign l_39[2325]    = ( l_40 [3349]);
assign l_39[2326]    = ( l_40 [3350]);
assign l_39[2327]    = ( l_40 [3351]);
assign l_39[2328]    = ( l_40 [3352]);
assign l_39[2329]    = ( l_40 [3353]);
assign l_39[2330]    = ( l_40 [3354]);
assign l_39[2331]    = ( l_40 [3355]);
assign l_39[2332]    = ( l_40 [3356]);
assign l_39[2333]    = ( l_40 [3357]);
assign l_39[2334]    = ( l_40 [3358]);
assign l_39[2335]    = ( l_40 [3359]);
assign l_39[2336]    = ( l_40 [3360]);
assign l_39[2337]    = ( l_40 [3361]);
assign l_39[2338]    = ( l_40 [3362]);
assign l_39[2339]    = ( l_40 [3363]);
assign l_39[2340]    = ( l_40 [3364]);
assign l_39[2341]    = ( l_40 [3365]);
assign l_39[2342]    = ( l_40 [3366]);
assign l_39[2343]    = ( l_40 [3367]);
assign l_39[2344]    = ( l_40 [3368]);
assign l_39[2345]    = ( l_40 [3369]);
assign l_39[2346]    = ( l_40 [3370]);
assign l_39[2347]    = ( l_40 [3371]);
assign l_39[2348]    = ( l_40 [3372]);
assign l_39[2349]    = ( l_40 [3373]);
assign l_39[2350]    = ( l_40 [3374]);
assign l_39[2351]    = ( l_40 [3375]);
assign l_39[2352]    = ( l_40 [3376]);
assign l_39[2353]    = ( l_40 [3377]);
assign l_39[2354]    = ( l_40 [3378]);
assign l_39[2355]    = ( l_40 [3379]);
assign l_39[2356]    = ( l_40 [3380]);
assign l_39[2357]    = ( l_40 [3381]);
assign l_39[2358]    = ( l_40 [3382]);
assign l_39[2359]    = ( l_40 [3383]);
assign l_39[2360]    = ( l_40 [3384]);
assign l_39[2361]    = ( l_40 [3385]);
assign l_39[2362]    = ( l_40 [3386]);
assign l_39[2363]    = ( l_40 [3387]);
assign l_39[2364]    = ( l_40 [3388]);
assign l_39[2365]    = ( l_40 [3389]);
assign l_39[2366]    = ( l_40 [3390]);
assign l_39[2367]    = ( l_40 [3391]);
assign l_39[2368]    = ( l_40 [3392]);
assign l_39[2369]    = ( l_40 [3393]);
assign l_39[2370]    = ( l_40 [3394]);
assign l_39[2371]    = ( l_40 [3395]);
assign l_39[2372]    = ( l_40 [3396]);
assign l_39[2373]    = ( l_40 [3397]);
assign l_39[2374]    = ( l_40 [3398]);
assign l_39[2375]    = ( l_40 [3399]);
assign l_39[2376]    = ( l_40 [3400]);
assign l_39[2377]    = ( l_40 [3401]);
assign l_39[2378]    = ( l_40 [3402]);
assign l_39[2379]    = ( l_40 [3403]);
assign l_39[2380]    = ( l_40 [3404]);
assign l_39[2381]    = ( l_40 [3405]);
assign l_39[2382]    = ( l_40 [3406]);
assign l_39[2383]    = ( l_40 [3407]);
assign l_39[2384]    = ( l_40 [3408]);
assign l_39[2385]    = ( l_40 [3409]);
assign l_39[2386]    = ( l_40 [3410]);
assign l_39[2387]    = ( l_40 [3411]);
assign l_39[2388]    = ( l_40 [3412]);
assign l_39[2389]    = ( l_40 [3413]);
assign l_39[2390]    = ( l_40 [3414]);
assign l_39[2391]    = ( l_40 [3415]);
assign l_39[2392]    = ( l_40 [3416]);
assign l_39[2393]    = ( l_40 [3417]);
assign l_39[2394]    = ( l_40 [3418]);
assign l_39[2395]    = ( l_40 [3419]);
assign l_39[2396]    = ( l_40 [3420]);
assign l_39[2397]    = ( l_40 [3421]);
assign l_39[2398]    = ( l_40 [3422]);
assign l_39[2399]    = ( l_40 [3423]);
assign l_39[2400]    = ( l_40 [3424]);
assign l_39[2401]    = ( l_40 [3425]);
assign l_39[2402]    = ( l_40 [3426]);
assign l_39[2403]    = ( l_40 [3427]);
assign l_39[2404]    = ( l_40 [3428]);
assign l_39[2405]    = ( l_40 [3429]);
assign l_39[2406]    = ( l_40 [3430]);
assign l_39[2407]    = ( l_40 [3431]);
assign l_39[2408]    = ( l_40 [3432]);
assign l_39[2409]    = ( l_40 [3433]);
assign l_39[2410]    = ( l_40 [3434]);
assign l_39[2411]    = ( l_40 [3435]);
assign l_39[2412]    = ( l_40 [3436]);
assign l_39[2413]    = ( l_40 [3437]);
assign l_39[2414]    = ( l_40 [3438]);
assign l_39[2415]    = ( l_40 [3439]);
assign l_39[2416]    = ( l_40 [3440]);
assign l_39[2417]    = ( l_40 [3441]);
assign l_39[2418]    = ( l_40 [3442]);
assign l_39[2419]    = ( l_40 [3443]);
assign l_39[2420]    = ( l_40 [3444]);
assign l_39[2421]    = ( l_40 [3445]);
assign l_39[2422]    = ( l_40 [3446]);
assign l_39[2423]    = ( l_40 [3447]);
assign l_39[2424]    = ( l_40 [3448]);
assign l_39[2425]    = ( l_40 [3449]);
assign l_39[2426]    = ( l_40 [3450]);
assign l_39[2427]    = ( l_40 [3451]);
assign l_39[2428]    = ( l_40 [3452]);
assign l_39[2429]    = ( l_40 [3453]);
assign l_39[2430]    = ( l_40 [3454]);
assign l_39[2431]    = ( l_40 [3455]);
assign l_39[2432]    = ( l_40 [3456]);
assign l_39[2433]    = ( l_40 [3457]);
assign l_39[2434]    = ( l_40 [3458]);
assign l_39[2435]    = ( l_40 [3459]);
assign l_39[2436]    = ( l_40 [3460]);
assign l_39[2437]    = ( l_40 [3461]);
assign l_39[2438]    = ( l_40 [3462]);
assign l_39[2439]    = ( l_40 [3463]);
assign l_39[2440]    = ( l_40 [3464]);
assign l_39[2441]    = ( l_40 [3465]);
assign l_39[2442]    = ( l_40 [3466]);
assign l_39[2443]    = ( l_40 [3467]);
assign l_39[2444]    = ( l_40 [3468]);
assign l_39[2445]    = ( l_40 [3469]);
assign l_39[2446]    = ( l_40 [3470]);
assign l_39[2447]    = ( l_40 [3471]);
assign l_39[2448]    = ( l_40 [3472]);
assign l_39[2449]    = ( l_40 [3473]);
assign l_39[2450]    = ( l_40 [3474]);
assign l_39[2451]    = ( l_40 [3475]);
assign l_39[2452]    = ( l_40 [3476]);
assign l_39[2453]    = ( l_40 [3477]);
assign l_39[2454]    = ( l_40 [3478]);
assign l_39[2455]    = ( l_40 [3479]);
assign l_39[2456]    = ( l_40 [3480]);
assign l_39[2457]    = ( l_40 [3481]);
assign l_39[2458]    = ( l_40 [3482]);
assign l_39[2459]    = ( l_40 [3483]);
assign l_39[2460]    = ( l_40 [3484]);
assign l_39[2461]    = ( l_40 [3485]);
assign l_39[2462]    = ( l_40 [3486]);
assign l_39[2463]    = ( l_40 [3487]);
assign l_39[2464]    = ( l_40 [3488]);
assign l_39[2465]    = ( l_40 [3489]);
assign l_39[2466]    = ( l_40 [3490]);
assign l_39[2467]    = ( l_40 [3491]);
assign l_39[2468]    = ( l_40 [3492]);
assign l_39[2469]    = ( l_40 [3493]);
assign l_39[2470]    = ( l_40 [3494]);
assign l_39[2471]    = ( l_40 [3495]);
assign l_39[2472]    = ( l_40 [3496]);
assign l_39[2473]    = ( l_40 [3497]);
assign l_39[2474]    = ( l_40 [3498]);
assign l_39[2475]    = ( l_40 [3499]);
assign l_39[2476]    = ( l_40 [3500]);
assign l_39[2477]    = ( l_40 [3501]);
assign l_39[2478]    = ( l_40 [3502]);
assign l_39[2479]    = ( l_40 [3503]);
assign l_39[2480]    = ( l_40 [3504]);
assign l_39[2481]    = ( l_40 [3505]);
assign l_39[2482]    = ( l_40 [3506]);
assign l_39[2483]    = ( l_40 [3507]);
assign l_39[2484]    = ( l_40 [3508]);
assign l_39[2485]    = ( l_40 [3509]);
assign l_39[2486]    = ( l_40 [3510]);
assign l_39[2487]    = ( l_40 [3511]);
assign l_39[2488]    = ( l_40 [3512]);
assign l_39[2489]    = ( l_40 [3513]);
assign l_39[2490]    = ( l_40 [3514]);
assign l_39[2491]    = ( l_40 [3515]);
assign l_39[2492]    = ( l_40 [3516]);
assign l_39[2493]    = ( l_40 [3517]);
assign l_39[2494]    = ( l_40 [3518]);
assign l_39[2495]    = ( l_40 [3519]);
assign l_39[2496]    = ( l_40 [3520]);
assign l_39[2497]    = ( l_40 [3521]);
assign l_39[2498]    = ( l_40 [3522]);
assign l_39[2499]    = ( l_40 [3523]);
assign l_39[2500]    = ( l_40 [3524]);
assign l_39[2501]    = ( l_40 [3525]);
assign l_39[2502]    = ( l_40 [3526]);
assign l_39[2503]    = ( l_40 [3527]);
assign l_39[2504]    = ( l_40 [3528]);
assign l_39[2505]    = ( l_40 [3529]);
assign l_39[2506]    = ( l_40 [3530]);
assign l_39[2507]    = ( l_40 [3531]);
assign l_39[2508]    = ( l_40 [3532]);
assign l_39[2509]    = ( l_40 [3533]);
assign l_39[2510]    = ( l_40 [3534]);
assign l_39[2511]    = ( l_40 [3535]);
assign l_39[2512]    = ( l_40 [3536]);
assign l_39[2513]    = ( l_40 [3537]);
assign l_39[2514]    = ( l_40 [3538]);
assign l_39[2515]    = ( l_40 [3539]);
assign l_39[2516]    = ( l_40 [3540]);
assign l_39[2517]    = ( l_40 [3541]);
assign l_39[2518]    = ( l_40 [3542]);
assign l_39[2519]    = ( l_40 [3543]);
assign l_39[2520]    = ( l_40 [3544]);
assign l_39[2521]    = ( l_40 [3545]);
assign l_39[2522]    = ( l_40 [3546]);
assign l_39[2523]    = ( l_40 [3547]);
assign l_39[2524]    = ( l_40 [3548]);
assign l_39[2525]    = ( l_40 [3549]);
assign l_39[2526]    = ( l_40 [3550]);
assign l_39[2527]    = ( l_40 [3551]);
assign l_39[2528]    = ( l_40 [3552]);
assign l_39[2529]    = ( l_40 [3553]);
assign l_39[2530]    = ( l_40 [3554]);
assign l_39[2531]    = ( l_40 [3555]);
assign l_39[2532]    = ( l_40 [3556]);
assign l_39[2533]    = ( l_40 [3557]);
assign l_39[2534]    = ( l_40 [3558]);
assign l_39[2535]    = ( l_40 [3559]);
assign l_39[2536]    = ( l_40 [3560]);
assign l_39[2537]    = ( l_40 [3561]);
assign l_39[2538]    = ( l_40 [3562]);
assign l_39[2539]    = ( l_40 [3563]);
assign l_39[2540]    = ( l_40 [3564]);
assign l_39[2541]    = ( l_40 [3565]);
assign l_39[2542]    = ( l_40 [3566]);
assign l_39[2543]    = ( l_40 [3567]);
assign l_39[2544]    = ( l_40 [3568]);
assign l_39[2545]    = ( l_40 [3569]);
assign l_39[2546]    = ( l_40 [3570]);
assign l_39[2547]    = ( l_40 [3571]);
assign l_39[2548]    = ( l_40 [3572]);
assign l_39[2549]    = ( l_40 [3573]);
assign l_39[2550]    = ( l_40 [3574]);
assign l_39[2551]    = ( l_40 [3575]);
assign l_39[2552]    = ( l_40 [3576]);
assign l_39[2553]    = ( l_40 [3577]);
assign l_39[2554]    = ( l_40 [3578]);
assign l_39[2555]    = ( l_40 [3579]);
assign l_39[2556]    = ( l_40 [3580]);
assign l_39[2557]    = ( l_40 [3581]);
assign l_39[2558]    = ( l_40 [3582]);
assign l_39[2559]    = ( l_40 [3583]);
assign l_39[2560]    = ( l_40 [3584]);
assign l_39[2561]    = ( l_40 [3585]);
assign l_39[2562]    = ( l_40 [3586]);
assign l_39[2563]    = ( l_40 [3587]);
assign l_39[2564]    = ( l_40 [3588]);
assign l_39[2565]    = ( l_40 [3589]);
assign l_39[2566]    = ( l_40 [3590]);
assign l_39[2567]    = ( l_40 [3591]);
assign l_39[2568]    = ( l_40 [3592]);
assign l_39[2569]    = ( l_40 [3593]);
assign l_39[2570]    = ( l_40 [3594]);
assign l_39[2571]    = ( l_40 [3595]);
assign l_39[2572]    = ( l_40 [3596]);
assign l_39[2573]    = ( l_40 [3597]);
assign l_39[2574]    = ( l_40 [3598]);
assign l_39[2575]    = ( l_40 [3599]);
assign l_39[2576]    = ( l_40 [3600]);
assign l_39[2577]    = ( l_40 [3601]);
assign l_39[2578]    = ( l_40 [3602]);
assign l_39[2579]    = ( l_40 [3603]);
assign l_39[2580]    = ( l_40 [3604]);
assign l_39[2581]    = ( l_40 [3605]);
assign l_39[2582]    = ( l_40 [3606]);
assign l_39[2583]    = ( l_40 [3607]);
assign l_39[2584]    = ( l_40 [3608]);
assign l_39[2585]    = ( l_40 [3609]);
assign l_39[2586]    = ( l_40 [3610]);
assign l_39[2587]    = ( l_40 [3611]);
assign l_39[2588]    = ( l_40 [3612]);
assign l_39[2589]    = ( l_40 [3613]);
assign l_39[2590]    = ( l_40 [3614]);
assign l_39[2591]    = ( l_40 [3615]);
assign l_39[2592]    = ( l_40 [3616]);
assign l_39[2593]    = ( l_40 [3617]);
assign l_39[2594]    = ( l_40 [3618]);
assign l_39[2595]    = ( l_40 [3619]);
assign l_39[2596]    = ( l_40 [3620]);
assign l_39[2597]    = ( l_40 [3621]);
assign l_39[2598]    = ( l_40 [3622]);
assign l_39[2599]    = ( l_40 [3623]);
assign l_39[2600]    = ( l_40 [3624]);
assign l_39[2601]    = ( l_40 [3625]);
assign l_39[2602]    = ( l_40 [3626]);
assign l_39[2603]    = ( l_40 [3627]);
assign l_39[2604]    = ( l_40 [3628]);
assign l_39[2605]    = ( l_40 [3629]);
assign l_39[2606]    = ( l_40 [3630]);
assign l_39[2607]    = ( l_40 [3631]);
assign l_39[2608]    = ( l_40 [3632]);
assign l_39[2609]    = ( l_40 [3633]);
assign l_39[2610]    = ( l_40 [3634]);
assign l_39[2611]    = ( l_40 [3635]);
assign l_39[2612]    = ( l_40 [3636]);
assign l_39[2613]    = ( l_40 [3637]);
assign l_39[2614]    = ( l_40 [3638]);
assign l_39[2615]    = ( l_40 [3639]);
assign l_39[2616]    = ( l_40 [3640]);
assign l_39[2617]    = ( l_40 [3641]);
assign l_39[2618]    = ( l_40 [3642]);
assign l_39[2619]    = ( l_40 [3643]);
assign l_39[2620]    = ( l_40 [3644]);
assign l_39[2621]    = ( l_40 [3645]);
assign l_39[2622]    = ( l_40 [3646]);
assign l_39[2623]    = ( l_40 [3647]);
assign l_39[2624]    = ( l_40 [3648]);
assign l_39[2625]    = ( l_40 [3649]);
assign l_39[2626]    = ( l_40 [3650]);
assign l_39[2627]    = ( l_40 [3651]);
assign l_39[2628]    = ( l_40 [3652]);
assign l_39[2629]    = ( l_40 [3653]);
assign l_39[2630]    = ( l_40 [3654]);
assign l_39[2631]    = ( l_40 [3655]);
assign l_39[2632]    = ( l_40 [3656]);
assign l_39[2633]    = ( l_40 [3657]);
assign l_39[2634]    = ( l_40 [3658]);
assign l_39[2635]    = ( l_40 [3659]);
assign l_39[2636]    = ( l_40 [3660]);
assign l_39[2637]    = ( l_40 [3661]);
assign l_39[2638]    = ( l_40 [3662]);
assign l_39[2639]    = ( l_40 [3663]);
assign l_39[2640]    = ( l_40 [3664]);
assign l_39[2641]    = ( l_40 [3665]);
assign l_39[2642]    = ( l_40 [3666]);
assign l_39[2643]    = ( l_40 [3667]);
assign l_39[2644]    = ( l_40 [3668]);
assign l_39[2645]    = ( l_40 [3669]);
assign l_39[2646]    = ( l_40 [3670]);
assign l_39[2647]    = ( l_40 [3671]);
assign l_39[2648]    = ( l_40 [3672]);
assign l_39[2649]    = ( l_40 [3673]);
assign l_39[2650]    = ( l_40 [3674]);
assign l_39[2651]    = ( l_40 [3675]);
assign l_39[2652]    = ( l_40 [3676]);
assign l_39[2653]    = ( l_40 [3677]);
assign l_39[2654]    = ( l_40 [3678]);
assign l_39[2655]    = ( l_40 [3679]);
assign l_39[2656]    = ( l_40 [3680]);
assign l_39[2657]    = ( l_40 [3681]);
assign l_39[2658]    = ( l_40 [3682]);
assign l_39[2659]    = ( l_40 [3683]);
assign l_39[2660]    = ( l_40 [3684]);
assign l_39[2661]    = ( l_40 [3685]);
assign l_39[2662]    = ( l_40 [3686]);
assign l_39[2663]    = ( l_40 [3687]);
assign l_39[2664]    = ( l_40 [3688]);
assign l_39[2665]    = ( l_40 [3689]);
assign l_39[2666]    = ( l_40 [3690]);
assign l_39[2667]    = ( l_40 [3691]);
assign l_39[2668]    = ( l_40 [3692]);
assign l_39[2669]    = ( l_40 [3693]);
assign l_39[2670]    = ( l_40 [3694]);
assign l_39[2671]    = ( l_40 [3695]);
assign l_39[2672]    = ( l_40 [3696]);
assign l_39[2673]    = ( l_40 [3697]);
assign l_39[2674]    = ( l_40 [3698]);
assign l_39[2675]    = ( l_40 [3699]);
assign l_39[2676]    = ( l_40 [3700]);
assign l_39[2677]    = ( l_40 [3701]);
assign l_39[2678]    = ( l_40 [3702]);
assign l_39[2679]    = ( l_40 [3703]);
assign l_39[2680]    = ( l_40 [3704]);
assign l_39[2681]    = ( l_40 [3705]);
assign l_39[2682]    = ( l_40 [3706]);
assign l_39[2683]    = ( l_40 [3707]);
assign l_39[2684]    = ( l_40 [3708]);
assign l_39[2685]    = ( l_40 [3709]);
assign l_39[2686]    = ( l_40 [3710]);
assign l_39[2687]    = ( l_40 [3711]);
assign l_39[2688]    = ( l_40 [3712]);
assign l_39[2689]    = ( l_40 [3713]);
assign l_39[2690]    = ( l_40 [3714]);
assign l_39[2691]    = ( l_40 [3715]);
assign l_39[2692]    = ( l_40 [3716]);
assign l_39[2693]    = ( l_40 [3717]);
assign l_39[2694]    = ( l_40 [3718]);
assign l_39[2695]    = ( l_40 [3719]);
assign l_39[2696]    = ( l_40 [3720]);
assign l_39[2697]    = ( l_40 [3721]);
assign l_39[2698]    = ( l_40 [3722]);
assign l_39[2699]    = ( l_40 [3723]);
assign l_39[2700]    = ( l_40 [3724]);
assign l_39[2701]    = ( l_40 [3725]);
assign l_39[2702]    = ( l_40 [3726]);
assign l_39[2703]    = ( l_40 [3727]);
assign l_39[2704]    = ( l_40 [3728]);
assign l_39[2705]    = ( l_40 [3729]);
assign l_39[2706]    = ( l_40 [3730]);
assign l_39[2707]    = ( l_40 [3731]);
assign l_39[2708]    = ( l_40 [3732]);
assign l_39[2709]    = ( l_40 [3733]);
assign l_39[2710]    = ( l_40 [3734]);
assign l_39[2711]    = ( l_40 [3735]);
assign l_39[2712]    = ( l_40 [3736]);
assign l_39[2713]    = ( l_40 [3737]);
assign l_39[2714]    = ( l_40 [3738]);
assign l_39[2715]    = ( l_40 [3739]);
assign l_39[2716]    = ( l_40 [3740]);
assign l_39[2717]    = ( l_40 [3741]);
assign l_39[2718]    = ( l_40 [3742]);
assign l_39[2719]    = ( l_40 [3743]);
assign l_39[2720]    = ( l_40 [3744]);
assign l_39[2721]    = ( l_40 [3745]);
assign l_39[2722]    = ( l_40 [3746]);
assign l_39[2723]    = ( l_40 [3747]);
assign l_39[2724]    = ( l_40 [3748]);
assign l_39[2725]    = ( l_40 [3749]);
assign l_39[2726]    = ( l_40 [3750]);
assign l_39[2727]    = ( l_40 [3751]);
assign l_39[2728]    = ( l_40 [3752]);
assign l_39[2729]    = ( l_40 [3753]);
assign l_39[2730]    = ( l_40 [3754]);
assign l_39[2731]    = ( l_40 [3755]);
assign l_39[2732]    = ( l_40 [3756]);
assign l_39[2733]    = ( l_40 [3757]);
assign l_39[2734]    = ( l_40 [3758]);
assign l_39[2735]    = ( l_40 [3759]);
assign l_39[2736]    = ( l_40 [3760]);
assign l_39[2737]    = ( l_40 [3761]);
assign l_39[2738]    = ( l_40 [3762]);
assign l_39[2739]    = ( l_40 [3763]);
assign l_39[2740]    = ( l_40 [3764]);
assign l_39[2741]    = ( l_40 [3765]);
assign l_39[2742]    = ( l_40 [3766]);
assign l_39[2743]    = ( l_40 [3767]);
assign l_39[2744]    = ( l_40 [3768]);
assign l_39[2745]    = ( l_40 [3769]);
assign l_39[2746]    = ( l_40 [3770]);
assign l_39[2747]    = ( l_40 [3771]);
assign l_39[2748]    = ( l_40 [3772]);
assign l_39[2749]    = ( l_40 [3773]);
assign l_39[2750]    = ( l_40 [3774]);
assign l_39[2751]    = ( l_40 [3775]);
assign l_39[2752]    = ( l_40 [3776]);
assign l_39[2753]    = ( l_40 [3777]);
assign l_39[2754]    = ( l_40 [3778]);
assign l_39[2755]    = ( l_40 [3779]);
assign l_39[2756]    = ( l_40 [3780]);
assign l_39[2757]    = ( l_40 [3781]);
assign l_39[2758]    = ( l_40 [3782]);
assign l_39[2759]    = ( l_40 [3783]);
assign l_39[2760]    = ( l_40 [3784]);
assign l_39[2761]    = ( l_40 [3785]);
assign l_39[2762]    = ( l_40 [3786]);
assign l_39[2763]    = ( l_40 [3787]);
assign l_39[2764]    = ( l_40 [3788]);
assign l_39[2765]    = ( l_40 [3789]);
assign l_39[2766]    = ( l_40 [3790]);
assign l_39[2767]    = ( l_40 [3791]);
assign l_39[2768]    = ( l_40 [3792]);
assign l_39[2769]    = ( l_40 [3793]);
assign l_39[2770]    = ( l_40 [3794]);
assign l_39[2771]    = ( l_40 [3795]);
assign l_39[2772]    = ( l_40 [3796]);
assign l_39[2773]    = ( l_40 [3797]);
assign l_39[2774]    = ( l_40 [3798]);
assign l_39[2775]    = ( l_40 [3799]);
assign l_39[2776]    = ( l_40 [3800]);
assign l_39[2777]    = ( l_40 [3801]);
assign l_39[2778]    = ( l_40 [3802]);
assign l_39[2779]    = ( l_40 [3803]);
assign l_39[2780]    = ( l_40 [3804]);
assign l_39[2781]    = ( l_40 [3805]);
assign l_39[2782]    = ( l_40 [3806]);
assign l_39[2783]    = ( l_40 [3807]);
assign l_39[2784]    = ( l_40 [3808]);
assign l_39[2785]    = ( l_40 [3809]);
assign l_39[2786]    = ( l_40 [3810]);
assign l_39[2787]    = ( l_40 [3811]);
assign l_39[2788]    = ( l_40 [3812]);
assign l_39[2789]    = ( l_40 [3813]);
assign l_39[2790]    = ( l_40 [3814]);
assign l_39[2791]    = ( l_40 [3815]);
assign l_39[2792]    = ( l_40 [3816]);
assign l_39[2793]    = ( l_40 [3817]);
assign l_39[2794]    = ( l_40 [3818]);
assign l_39[2795]    = ( l_40 [3819]);
assign l_39[2796]    = ( l_40 [3820]);
assign l_39[2797]    = ( l_40 [3821]);
assign l_39[2798]    = ( l_40 [3822]);
assign l_39[2799]    = ( l_40 [3823]);
assign l_39[2800]    = ( l_40 [3824]);
assign l_39[2801]    = ( l_40 [3825]);
assign l_39[2802]    = ( l_40 [3826]);
assign l_39[2803]    = ( l_40 [3827]);
assign l_39[2804]    = ( l_40 [3828]);
assign l_39[2805]    = ( l_40 [3829]);
assign l_39[2806]    = ( l_40 [3830]);
assign l_39[2807]    = ( l_40 [3831]);
assign l_39[2808]    = ( l_40 [3832]);
assign l_39[2809]    = ( l_40 [3833]);
assign l_39[2810]    = ( l_40 [3834]);
assign l_39[2811]    = ( l_40 [3835]);
assign l_39[2812]    = ( l_40 [3836]);
assign l_39[2813]    = ( l_40 [3837]);
assign l_39[2814]    = ( l_40 [3838]);
assign l_39[2815]    = ( l_40 [3839]);
assign l_39[2816]    = ( l_40 [3840]);
assign l_39[2817]    = ( l_40 [3841]);
assign l_39[2818]    = ( l_40 [3842]);
assign l_39[2819]    = ( l_40 [3843]);
assign l_39[2820]    = ( l_40 [3844]);
assign l_39[2821]    = ( l_40 [3845]);
assign l_39[2822]    = ( l_40 [3846]);
assign l_39[2823]    = ( l_40 [3847]);
assign l_39[2824]    = ( l_40 [3848]);
assign l_39[2825]    = ( l_40 [3849]);
assign l_39[2826]    = ( l_40 [3850]);
assign l_39[2827]    = ( l_40 [3851]);
assign l_39[2828]    = ( l_40 [3852]);
assign l_39[2829]    = ( l_40 [3853]);
assign l_39[2830]    = ( l_40 [3854]);
assign l_39[2831]    = ( l_40 [3855]);
assign l_39[2832]    = ( l_40 [3856]);
assign l_39[2833]    = ( l_40 [3857]);
assign l_39[2834]    = ( l_40 [3858]);
assign l_39[2835]    = ( l_40 [3859]);
assign l_39[2836]    = ( l_40 [3860]);
assign l_39[2837]    = ( l_40 [3861]);
assign l_39[2838]    = ( l_40 [3862]);
assign l_39[2839]    = ( l_40 [3863]);
assign l_39[2840]    = ( l_40 [3864]);
assign l_39[2841]    = ( l_40 [3865]);
assign l_39[2842]    = ( l_40 [3866]);
assign l_39[2843]    = ( l_40 [3867]);
assign l_39[2844]    = ( l_40 [3868]);
assign l_39[2845]    = ( l_40 [3869]);
assign l_39[2846]    = ( l_40 [3870]);
assign l_39[2847]    = ( l_40 [3871]);
assign l_39[2848]    = ( l_40 [3872]);
assign l_39[2849]    = ( l_40 [3873]);
assign l_39[2850]    = ( l_40 [3874]);
assign l_39[2851]    = ( l_40 [3875]);
assign l_39[2852]    = ( l_40 [3876]);
assign l_39[2853]    = ( l_40 [3877]);
assign l_39[2854]    = ( l_40 [3878]);
assign l_39[2855]    = ( l_40 [3879]);
assign l_39[2856]    = ( l_40 [3880]);
assign l_39[2857]    = ( l_40 [3881]);
assign l_39[2858]    = ( l_40 [3882]);
assign l_39[2859]    = ( l_40 [3883]);
assign l_39[2860]    = ( l_40 [3884]);
assign l_39[2861]    = ( l_40 [3885]);
assign l_39[2862]    = ( l_40 [3886]);
assign l_39[2863]    = ( l_40 [3887]);
assign l_39[2864]    = ( l_40 [3888]);
assign l_39[2865]    = ( l_40 [3889]);
assign l_39[2866]    = ( l_40 [3890]);
assign l_39[2867]    = ( l_40 [3891]);
assign l_39[2868]    = ( l_40 [3892]);
assign l_39[2869]    = ( l_40 [3893]);
assign l_39[2870]    = ( l_40 [3894]);
assign l_39[2871]    = ( l_40 [3895]);
assign l_39[2872]    = ( l_40 [3896]);
assign l_39[2873]    = ( l_40 [3897]);
assign l_39[2874]    = ( l_40 [3898]);
assign l_39[2875]    = ( l_40 [3899]);
assign l_39[2876]    = ( l_40 [3900]);
assign l_39[2877]    = ( l_40 [3901]);
assign l_39[2878]    = ( l_40 [3902]);
assign l_39[2879]    = ( l_40 [3903]);
assign l_39[2880]    = ( l_40 [3904]);
assign l_39[2881]    = ( l_40 [3905]);
assign l_39[2882]    = ( l_40 [3906]);
assign l_39[2883]    = ( l_40 [3907]);
assign l_39[2884]    = ( l_40 [3908]);
assign l_39[2885]    = ( l_40 [3909]);
assign l_39[2886]    = ( l_40 [3910]);
assign l_39[2887]    = ( l_40 [3911]);
assign l_39[2888]    = ( l_40 [3912]);
assign l_39[2889]    = ( l_40 [3913]);
assign l_39[2890]    = ( l_40 [3914]);
assign l_39[2891]    = ( l_40 [3915]);
assign l_39[2892]    = ( l_40 [3916]);
assign l_39[2893]    = ( l_40 [3917]);
assign l_39[2894]    = ( l_40 [3918]);
assign l_39[2895]    = ( l_40 [3919]);
assign l_39[2896]    = ( l_40 [3920]);
assign l_39[2897]    = ( l_40 [3921]);
assign l_39[2898]    = ( l_40 [3922]);
assign l_39[2899]    = ( l_40 [3923]);
assign l_39[2900]    = ( l_40 [3924]);
assign l_39[2901]    = ( l_40 [3925]);
assign l_39[2902]    = ( l_40 [3926]);
assign l_39[2903]    = ( l_40 [3927]);
assign l_39[2904]    = ( l_40 [3928]);
assign l_39[2905]    = ( l_40 [3929]);
assign l_39[2906]    = ( l_40 [3930]);
assign l_39[2907]    = ( l_40 [3931]);
assign l_39[2908]    = ( l_40 [3932]);
assign l_39[2909]    = ( l_40 [3933]);
assign l_39[2910]    = ( l_40 [3934]);
assign l_39[2911]    = ( l_40 [3935]);
assign l_39[2912]    = ( l_40 [3936]);
assign l_39[2913]    = ( l_40 [3937]);
assign l_39[2914]    = ( l_40 [3938]);
assign l_39[2915]    = ( l_40 [3939]);
assign l_39[2916]    = ( l_40 [3940]);
assign l_39[2917]    = ( l_40 [3941]);
assign l_39[2918]    = ( l_40 [3942]);
assign l_39[2919]    = ( l_40 [3943]);
assign l_39[2920]    = ( l_40 [3944]);
assign l_39[2921]    = ( l_40 [3945]);
assign l_39[2922]    = ( l_40 [3946]);
assign l_39[2923]    = ( l_40 [3947]);
assign l_39[2924]    = ( l_40 [3948]);
assign l_39[2925]    = ( l_40 [3949]);
assign l_39[2926]    = ( l_40 [3950]);
assign l_39[2927]    = ( l_40 [3951]);
assign l_39[2928]    = ( l_40 [3952]);
assign l_39[2929]    = ( l_40 [3953]);
assign l_39[2930]    = ( l_40 [3954]);
assign l_39[2931]    = ( l_40 [3955]);
assign l_39[2932]    = ( l_40 [3956]);
assign l_39[2933]    = ( l_40 [3957]);
assign l_39[2934]    = ( l_40 [3958]);
assign l_39[2935]    = ( l_40 [3959]);
assign l_39[2936]    = ( l_40 [3960]);
assign l_39[2937]    = ( l_40 [3961]);
assign l_39[2938]    = ( l_40 [3962]);
assign l_39[2939]    = ( l_40 [3963]);
assign l_39[2940]    = ( l_40 [3964]);
assign l_39[2941]    = ( l_40 [3965]);
assign l_39[2942]    = ( l_40 [3966]);
assign l_39[2943]    = ( l_40 [3967]);
assign l_39[2944]    = ( l_40 [3968]);
assign l_39[2945]    = ( l_40 [3969]);
assign l_39[2946]    = ( l_40 [3970]);
assign l_39[2947]    = ( l_40 [3971]);
assign l_39[2948]    = ( l_40 [3972]);
assign l_39[2949]    = ( l_40 [3973]);
assign l_39[2950]    = ( l_40 [3974]);
assign l_39[2951]    = ( l_40 [3975]);
assign l_39[2952]    = ( l_40 [3976]);
assign l_39[2953]    = ( l_40 [3977]);
assign l_39[2954]    = ( l_40 [3978]);
assign l_39[2955]    = ( l_40 [3979]);
assign l_39[2956]    = ( l_40 [3980]);
assign l_39[2957]    = ( l_40 [3981]);
assign l_39[2958]    = ( l_40 [3982]);
assign l_39[2959]    = ( l_40 [3983]);
assign l_39[2960]    = ( l_40 [3984]);
assign l_39[2961]    = ( l_40 [3985]);
assign l_39[2962]    = ( l_40 [3986]);
assign l_39[2963]    = ( l_40 [3987]);
assign l_39[2964]    = ( l_40 [3988]);
assign l_39[2965]    = ( l_40 [3989]);
assign l_39[2966]    = ( l_40 [3990]);
assign l_39[2967]    = ( l_40 [3991]);
assign l_39[2968]    = ( l_40 [3992]);
assign l_39[2969]    = ( l_40 [3993]);
assign l_39[2970]    = ( l_40 [3994]);
assign l_39[2971]    = ( l_40 [3995]);
assign l_39[2972]    = ( l_40 [3996]);
assign l_39[2973]    = ( l_40 [3997]);
assign l_39[2974]    = ( l_40 [3998]);
assign l_39[2975]    = ( l_40 [3999]);
assign l_39[2976]    = ( l_40 [4000]);
assign l_39[2977]    = ( l_40 [4001]);
assign l_39[2978]    = ( l_40 [4002]);
assign l_39[2979]    = ( l_40 [4003]);
assign l_39[2980]    = ( l_40 [4004]);
assign l_39[2981]    = ( l_40 [4005]);
assign l_39[2982]    = ( l_40 [4006]);
assign l_39[2983]    = ( l_40 [4007]);
assign l_39[2984]    = ( l_40 [4008]);
assign l_39[2985]    = ( l_40 [4009]);
assign l_39[2986]    = ( l_40 [4010]);
assign l_39[2987]    = ( l_40 [4011]);
assign l_39[2988]    = ( l_40 [4012]);
assign l_39[2989]    = ( l_40 [4013]);
assign l_39[2990]    = ( l_40 [4014]);
assign l_39[2991]    = ( l_40 [4015]);
assign l_39[2992]    = ( l_40 [4016]);
assign l_39[2993]    = ( l_40 [4017]);
assign l_39[2994]    = ( l_40 [4018]);
assign l_39[2995]    = ( l_40 [4019]);
assign l_39[2996]    = ( l_40 [4020]);
assign l_39[2997]    = ( l_40 [4021]);
assign l_39[2998]    = ( l_40 [4022]);
assign l_39[2999]    = ( l_40 [4023]);
assign l_39[3000]    = ( l_40 [4024]);
assign l_39[3001]    = ( l_40 [4025]);
assign l_39[3002]    = ( l_40 [4026]);
assign l_39[3003]    = ( l_40 [4027]);
assign l_39[3004]    = ( l_40 [4028]);
assign l_39[3005]    = ( l_40 [4029]);
assign l_39[3006]    = ( l_40 [4030]);
assign l_39[3007]    = ( l_40 [4031]);
assign l_39[3008]    = ( l_40 [4032]);
assign l_39[3009]    = ( l_40 [4033]);
assign l_39[3010]    = ( l_40 [4034]);
assign l_39[3011]    = ( l_40 [4035]);
assign l_39[3012]    = ( l_40 [4036]);
assign l_39[3013]    = ( l_40 [4037]);
assign l_39[3014]    = ( l_40 [4038]);
assign l_39[3015]    = ( l_40 [4039]);
assign l_39[3016]    = ( l_40 [4040]);
assign l_39[3017]    = ( l_40 [4041]);
assign l_39[3018]    = ( l_40 [4042]);
assign l_39[3019]    = ( l_40 [4043]);
assign l_39[3020]    = ( l_40 [4044]);
assign l_39[3021]    = ( l_40 [4045]);
assign l_39[3022]    = ( l_40 [4046]);
assign l_39[3023]    = ( l_40 [4047]);
assign l_39[3024]    = ( l_40 [4048]);
assign l_39[3025]    = ( l_40 [4049]);
assign l_39[3026]    = ( l_40 [4050]);
assign l_39[3027]    = ( l_40 [4051]);
assign l_39[3028]    = ( l_40 [4052]);
assign l_39[3029]    = ( l_40 [4053]);
assign l_39[3030]    = ( l_40 [4054]);
assign l_39[3031]    = ( l_40 [4055]);
assign l_39[3032]    = ( l_40 [4056]);
assign l_39[3033]    = ( l_40 [4057]);
assign l_39[3034]    = ( l_40 [4058]);
assign l_39[3035]    = ( l_40 [4059]);
assign l_39[3036]    = ( l_40 [4060]);
assign l_39[3037]    = ( l_40 [4061]);
assign l_39[3038]    = ( l_40 [4062]);
assign l_39[3039]    = ( l_40 [4063]);
assign l_39[3040]    = ( l_40 [4064]);
assign l_39[3041]    = ( l_40 [4065]);
assign l_39[3042]    = ( l_40 [4066]);
assign l_39[3043]    = ( l_40 [4067]);
assign l_39[3044]    = ( l_40 [4068]);
assign l_39[3045]    = ( l_40 [4069]);
assign l_39[3046]    = ( l_40 [4070]);
assign l_39[3047]    = ( l_40 [4071]);
assign l_39[3048]    = ( l_40 [4072]);
assign l_39[3049]    = ( l_40 [4073]);
assign l_39[3050]    = ( l_40 [4074]);
assign l_39[3051]    = ( l_40 [4075]);
assign l_39[3052]    = ( l_40 [4076]);
assign l_39[3053]    = ( l_40 [4077]);
assign l_39[3054]    = ( l_40 [4078]);
assign l_39[3055]    = ( l_40 [4079]);
assign l_39[3056]    = ( l_40 [4080]);
assign l_39[3057]    = ( l_40 [4081]);
assign l_39[3058]    = ( l_40 [4082]);
assign l_39[3059]    = ( l_40 [4083]);
assign l_39[3060]    = ( l_40 [4084]);
assign l_39[3061]    = ( l_40 [4085]);
assign l_39[3062]    = ( l_40 [4086]);
assign l_39[3063]    = ( l_40 [4087]);
assign l_39[3064]    = ( l_40 [4088]);
assign l_39[3065]    = ( l_40 [4089]);
assign l_39[3066]    = ( l_40 [4090]);
assign l_39[3067]    = ( l_40 [4091]);
assign l_39[3068]    = ( l_40 [4092]);
assign l_39[3069]    = ( l_40 [4093]);
assign l_39[3070]    = ( l_40 [4094]);
assign l_39[3071]    = ( l_40 [4095]);
assign l_39[3072]    = ( l_40 [4096]);
assign l_39[3073]    = ( l_40 [4097]);
assign l_39[3074]    = ( l_40 [4098]);
assign l_39[3075]    = ( l_40 [4099]);
assign l_39[3076]    = ( l_40 [4100]);
assign l_39[3077]    = ( l_40 [4101]);
assign l_39[3078]    = ( l_40 [4102]);
assign l_39[3079]    = ( l_40 [4103]);
assign l_39[3080]    = ( l_40 [4104]);
assign l_39[3081]    = ( l_40 [4105]);
assign l_39[3082]    = ( l_40 [4106]);
assign l_39[3083]    = ( l_40 [4107]);
assign l_39[3084]    = ( l_40 [4108]);
assign l_39[3085]    = ( l_40 [4109]);
assign l_39[3086]    = ( l_40 [4110]);
assign l_39[3087]    = ( l_40 [4111]);
assign l_39[3088]    = ( l_40 [4112]);
assign l_39[3089]    = ( l_40 [4113]);
assign l_40[0]    = ( l_41 [0]);
assign l_40[1]    = ( l_41 [1] & !i[1819]) | ( l_41 [2] &  i[1819]);
assign l_40[2]    = ( l_41 [3] & !i[1819]) | ( l_41 [4] &  i[1819]);
assign l_40[3]    = ( l_41 [5] & !i[1819]) | ( l_41 [6] &  i[1819]);
assign l_40[4]    = ( l_41 [7] & !i[1819]) | ( l_41 [8] &  i[1819]);
assign l_40[5]    = ( l_41 [9] & !i[1819]) | ( l_41 [10] &  i[1819]);
assign l_40[6]    = ( l_41 [11] & !i[1819]) | ( l_41 [12] &  i[1819]);
assign l_40[7]    = ( l_41 [13] & !i[1819]) | ( l_41 [14] &  i[1819]);
assign l_40[8]    = ( l_41 [15] & !i[1819]) | ( l_41 [16] &  i[1819]);
assign l_40[9]    = ( l_41 [17] & !i[1819]) | ( l_41 [18] &  i[1819]);
assign l_40[10]    = ( l_41 [19]);
assign l_40[11]    = ( l_41 [20] & !i[1819]) | ( l_41 [21] &  i[1819]);
assign l_40[12]    = ( l_41 [22] & !i[1819]) | ( l_41 [23] &  i[1819]);
assign l_40[13]    = ( l_41 [24] & !i[1819]) | ( l_41 [25] &  i[1819]);
assign l_40[14]    = ( l_41 [26] & !i[1819]) | ( l_41 [27] &  i[1819]);
assign l_40[15]    = ( l_41 [28] & !i[1819]) | ( l_41 [29] &  i[1819]);
assign l_40[16]    = ( l_41 [30] & !i[1819]) | ( l_41 [31] &  i[1819]);
assign l_40[17]    = ( l_41 [32] & !i[1819]) | ( l_41 [33] &  i[1819]);
assign l_40[18]    = ( l_41 [34] & !i[1819]) | ( l_41 [35] &  i[1819]);
assign l_40[19]    = ( l_41 [36] & !i[1819]) | ( l_41 [37] &  i[1819]);
assign l_40[20]    = ( l_41 [38] & !i[1819]) | ( l_41 [39] &  i[1819]);
assign l_40[21]    = ( l_41 [40] & !i[1819]) | ( l_41 [41] &  i[1819]);
assign l_40[22]    = ( l_41 [42] & !i[1819]) | ( l_41 [43] &  i[1819]);
assign l_40[23]    = ( l_41 [44] & !i[1819]) | ( l_41 [45] &  i[1819]);
assign l_40[24]    = ( l_41 [46] & !i[1819]) | ( l_41 [47] &  i[1819]);
assign l_40[25]    = ( l_41 [48] & !i[1819]) | ( l_41 [49] &  i[1819]);
assign l_40[26]    = ( l_41 [50] & !i[1819]) | ( l_41 [51] &  i[1819]);
assign l_40[27]    = ( l_41 [52] & !i[1819]) | ( l_41 [53] &  i[1819]);
assign l_40[28]    = ( l_41 [54] & !i[1819]) | ( l_41 [55] &  i[1819]);
assign l_40[29]    = ( l_41 [56] & !i[1819]) | ( l_41 [57] &  i[1819]);
assign l_40[30]    = ( l_41 [58] & !i[1819]) | ( l_41 [59] &  i[1819]);
assign l_40[31]    = ( l_41 [60] & !i[1819]) | ( l_41 [61] &  i[1819]);
assign l_40[32]    = ( l_41 [62] & !i[1819]) | ( l_41 [63] &  i[1819]);
assign l_40[33]    = ( l_41 [64] & !i[1819]) | ( l_41 [65] &  i[1819]);
assign l_40[34]    = ( l_41 [66] & !i[1819]) | ( l_41 [67] &  i[1819]);
assign l_40[35]    = ( l_41 [68] & !i[1819]) | ( l_41 [69] &  i[1819]);
assign l_40[36]    = ( l_41 [70] & !i[1819]) | ( l_41 [71] &  i[1819]);
assign l_40[37]    = ( l_41 [72] & !i[1819]) | ( l_41 [73] &  i[1819]);
assign l_40[38]    = ( l_41 [74] & !i[1819]) | ( l_41 [75] &  i[1819]);
assign l_40[39]    = ( l_41 [76] & !i[1819]) | ( l_41 [77] &  i[1819]);
assign l_40[40]    = ( l_41 [78] & !i[1819]) | ( l_41 [79] &  i[1819]);
assign l_40[41]    = ( l_41 [80] & !i[1819]) | ( l_41 [81] &  i[1819]);
assign l_40[42]    = ( l_41 [82] & !i[1819]) | ( l_41 [83] &  i[1819]);
assign l_40[43]    = ( l_41 [84] & !i[1819]) | ( l_41 [85] &  i[1819]);
assign l_40[44]    = ( l_41 [86] & !i[1819]) | ( l_41 [87] &  i[1819]);
assign l_40[45]    = ( l_41 [88] & !i[1819]) | ( l_41 [89] &  i[1819]);
assign l_40[46]    = ( l_41 [90] & !i[1819]) | ( l_41 [91] &  i[1819]);
assign l_40[47]    = ( l_41 [92] & !i[1819]) | ( l_41 [93] &  i[1819]);
assign l_40[48]    = ( l_41 [94] & !i[1819]) | ( l_41 [95] &  i[1819]);
assign l_40[49]    = ( l_41 [96] & !i[1819]) | ( l_41 [97] &  i[1819]);
assign l_40[50]    = ( l_41 [98] & !i[1819]) | ( l_41 [99] &  i[1819]);
assign l_40[51]    = ( l_41 [100] & !i[1819]) | ( l_41 [101] &  i[1819]);
assign l_40[52]    = ( l_41 [102] & !i[1819]) | ( l_41 [103] &  i[1819]);
assign l_40[53]    = ( l_41 [104] & !i[1819]) | ( l_41 [105] &  i[1819]);
assign l_40[54]    = ( l_41 [106] & !i[1819]) | ( l_41 [107] &  i[1819]);
assign l_40[55]    = ( l_41 [108] & !i[1819]) | ( l_41 [109] &  i[1819]);
assign l_40[56]    = ( l_41 [110] & !i[1819]) | ( l_41 [111] &  i[1819]);
assign l_40[57]    = ( l_41 [112] & !i[1819]) | ( l_41 [113] &  i[1819]);
assign l_40[58]    = ( l_41 [114] & !i[1819]) | ( l_41 [115] &  i[1819]);
assign l_40[59]    = ( l_41 [116] & !i[1819]) | ( l_41 [117] &  i[1819]);
assign l_40[60]    = ( l_41 [118] & !i[1819]) | ( l_41 [119] &  i[1819]);
assign l_40[61]    = ( l_41 [120] & !i[1819]) | ( l_41 [121] &  i[1819]);
assign l_40[62]    = ( l_41 [122] & !i[1819]) | ( l_41 [123] &  i[1819]);
assign l_40[63]    = ( l_41 [124] & !i[1819]) | ( l_41 [125] &  i[1819]);
assign l_40[64]    = ( l_41 [126] & !i[1819]) | ( l_41 [127] &  i[1819]);
assign l_40[65]    = ( l_41 [128] & !i[1819]) | ( l_41 [129] &  i[1819]);
assign l_40[66]    = ( l_41 [130] & !i[1819]) | ( l_41 [131] &  i[1819]);
assign l_40[67]    = ( l_41 [132] & !i[1819]) | ( l_41 [133] &  i[1819]);
assign l_40[68]    = ( l_41 [134] & !i[1819]) | ( l_41 [135] &  i[1819]);
assign l_40[69]    = ( l_41 [136] & !i[1819]) | ( l_41 [137] &  i[1819]);
assign l_40[70]    = ( l_41 [138] & !i[1819]) | ( l_41 [139] &  i[1819]);
assign l_40[71]    = ( l_41 [140] & !i[1819]) | ( l_41 [141] &  i[1819]);
assign l_40[72]    = ( l_41 [142] & !i[1819]) | ( l_41 [143] &  i[1819]);
assign l_40[73]    = ( l_41 [144] & !i[1819]) | ( l_41 [145] &  i[1819]);
assign l_40[74]    = ( l_41 [146] & !i[1819]) | ( l_41 [147] &  i[1819]);
assign l_40[75]    = ( l_41 [148] & !i[1819]) | ( l_41 [149] &  i[1819]);
assign l_40[76]    = ( l_41 [150] & !i[1819]) | ( l_41 [151] &  i[1819]);
assign l_40[77]    = ( l_41 [152] & !i[1819]) | ( l_41 [153] &  i[1819]);
assign l_40[78]    = ( l_41 [154] & !i[1819]) | ( l_41 [155] &  i[1819]);
assign l_40[79]    = ( l_41 [156] & !i[1819]) | ( l_41 [157] &  i[1819]);
assign l_40[80]    = ( l_41 [158] & !i[1819]) | ( l_41 [159] &  i[1819]);
assign l_40[81]    = ( l_41 [160] & !i[1819]) | ( l_41 [161] &  i[1819]);
assign l_40[82]    = ( l_41 [162] & !i[1819]) | ( l_41 [163] &  i[1819]);
assign l_40[83]    = ( l_41 [164] & !i[1819]) | ( l_41 [165] &  i[1819]);
assign l_40[84]    = ( l_41 [166] & !i[1819]) | ( l_41 [167] &  i[1819]);
assign l_40[85]    = ( l_41 [168] & !i[1819]) | ( l_41 [169] &  i[1819]);
assign l_40[86]    = ( l_41 [170] & !i[1819]) | ( l_41 [171] &  i[1819]);
assign l_40[87]    = ( l_41 [172] & !i[1819]) | ( l_41 [173] &  i[1819]);
assign l_40[88]    = ( l_41 [174] & !i[1819]) | ( l_41 [175] &  i[1819]);
assign l_40[89]    = ( l_41 [176] & !i[1819]) | ( l_41 [177] &  i[1819]);
assign l_40[90]    = ( l_41 [178] & !i[1819]) | ( l_41 [179] &  i[1819]);
assign l_40[91]    = ( l_41 [180] & !i[1819]) | ( l_41 [181] &  i[1819]);
assign l_40[92]    = ( l_41 [182] & !i[1819]) | ( l_41 [183] &  i[1819]);
assign l_40[93]    = ( l_41 [184] & !i[1819]) | ( l_41 [185] &  i[1819]);
assign l_40[94]    = ( l_41 [186] & !i[1819]) | ( l_41 [187] &  i[1819]);
assign l_40[95]    = ( l_41 [188] & !i[1819]) | ( l_41 [189] &  i[1819]);
assign l_40[96]    = ( l_41 [190] & !i[1819]) | ( l_41 [191] &  i[1819]);
assign l_40[97]    = ( l_41 [192] & !i[1819]) | ( l_41 [193] &  i[1819]);
assign l_40[98]    = ( l_41 [194] & !i[1819]) | ( l_41 [195] &  i[1819]);
assign l_40[99]    = ( l_41 [196] & !i[1819]) | ( l_41 [197] &  i[1819]);
assign l_40[100]    = ( l_41 [198] & !i[1819]) | ( l_41 [199] &  i[1819]);
assign l_40[101]    = ( l_41 [200] & !i[1819]) | ( l_41 [201] &  i[1819]);
assign l_40[102]    = ( l_41 [202] & !i[1819]) | ( l_41 [203] &  i[1819]);
assign l_40[103]    = ( l_41 [204] & !i[1819]) | ( l_41 [205] &  i[1819]);
assign l_40[104]    = ( l_41 [206] & !i[1819]) | ( l_41 [207] &  i[1819]);
assign l_40[105]    = ( l_41 [208] & !i[1819]) | ( l_41 [209] &  i[1819]);
assign l_40[106]    = ( l_41 [210] & !i[1819]) | ( l_41 [211] &  i[1819]);
assign l_40[107]    = ( l_41 [212] & !i[1819]) | ( l_41 [213] &  i[1819]);
assign l_40[108]    = ( l_41 [214] & !i[1819]) | ( l_41 [215] &  i[1819]);
assign l_40[109]    = ( l_41 [216] & !i[1819]) | ( l_41 [217] &  i[1819]);
assign l_40[110]    = ( l_41 [218] & !i[1819]) | ( l_41 [219] &  i[1819]);
assign l_40[111]    = ( l_41 [220] & !i[1819]) | ( l_41 [221] &  i[1819]);
assign l_40[112]    = ( l_41 [222] & !i[1819]) | ( l_41 [223] &  i[1819]);
assign l_40[113]    = ( l_41 [224] & !i[1819]) | ( l_41 [225] &  i[1819]);
assign l_40[114]    = ( l_41 [226] & !i[1819]) | ( l_41 [227] &  i[1819]);
assign l_40[115]    = ( l_41 [228] & !i[1819]) | ( l_41 [229] &  i[1819]);
assign l_40[116]    = ( l_41 [230] & !i[1819]) | ( l_41 [231] &  i[1819]);
assign l_40[117]    = ( l_41 [232] & !i[1819]) | ( l_41 [233] &  i[1819]);
assign l_40[118]    = ( l_41 [234] & !i[1819]) | ( l_41 [235] &  i[1819]);
assign l_40[119]    = ( l_41 [236] & !i[1819]) | ( l_41 [237] &  i[1819]);
assign l_40[120]    = ( l_41 [238] & !i[1819]) | ( l_41 [239] &  i[1819]);
assign l_40[121]    = ( l_41 [240] & !i[1819]) | ( l_41 [241] &  i[1819]);
assign l_40[122]    = ( l_41 [242] & !i[1819]) | ( l_41 [243] &  i[1819]);
assign l_40[123]    = ( l_41 [244] & !i[1819]) | ( l_41 [245] &  i[1819]);
assign l_40[124]    = ( l_41 [246] & !i[1819]) | ( l_41 [247] &  i[1819]);
assign l_40[125]    = ( l_41 [248] & !i[1819]) | ( l_41 [249] &  i[1819]);
assign l_40[126]    = ( l_41 [250] & !i[1819]) | ( l_41 [251] &  i[1819]);
assign l_40[127]    = ( l_41 [252] & !i[1819]) | ( l_41 [253] &  i[1819]);
assign l_40[128]    = ( l_41 [254] & !i[1819]) | ( l_41 [255] &  i[1819]);
assign l_40[129]    = ( l_41 [256] & !i[1819]) | ( l_41 [257] &  i[1819]);
assign l_40[130]    = ( l_41 [258] & !i[1819]) | ( l_41 [259] &  i[1819]);
assign l_40[131]    = ( l_41 [260] & !i[1819]) | ( l_41 [261] &  i[1819]);
assign l_40[132]    = ( l_41 [262] & !i[1819]) | ( l_41 [263] &  i[1819]);
assign l_40[133]    = ( l_41 [264] & !i[1819]) | ( l_41 [265] &  i[1819]);
assign l_40[134]    = ( l_41 [266] & !i[1819]) | ( l_41 [267] &  i[1819]);
assign l_40[135]    = ( l_41 [268] & !i[1819]) | ( l_41 [269] &  i[1819]);
assign l_40[136]    = ( l_41 [270] & !i[1819]) | ( l_41 [271] &  i[1819]);
assign l_40[137]    = ( l_41 [272] & !i[1819]) | ( l_41 [273] &  i[1819]);
assign l_40[138]    = ( l_41 [274] & !i[1819]) | ( l_41 [275] &  i[1819]);
assign l_40[139]    = ( l_41 [276] & !i[1819]) | ( l_41 [277] &  i[1819]);
assign l_40[140]    = ( l_41 [278] & !i[1819]) | ( l_41 [279] &  i[1819]);
assign l_40[141]    = ( l_41 [280] & !i[1819]) | ( l_41 [281] &  i[1819]);
assign l_40[142]    = ( l_41 [282] & !i[1819]) | ( l_41 [283] &  i[1819]);
assign l_40[143]    = ( l_41 [284] & !i[1819]) | ( l_41 [285] &  i[1819]);
assign l_40[144]    = ( l_41 [286] & !i[1819]) | ( l_41 [287] &  i[1819]);
assign l_40[145]    = ( l_41 [288] & !i[1819]) | ( l_41 [289] &  i[1819]);
assign l_40[146]    = ( l_41 [290] & !i[1819]) | ( l_41 [291] &  i[1819]);
assign l_40[147]    = ( l_41 [292] & !i[1819]) | ( l_41 [293] &  i[1819]);
assign l_40[148]    = ( l_41 [294] & !i[1819]) | ( l_41 [295] &  i[1819]);
assign l_40[149]    = ( l_41 [296] & !i[1819]) | ( l_41 [297] &  i[1819]);
assign l_40[150]    = ( l_41 [298] & !i[1819]) | ( l_41 [299] &  i[1819]);
assign l_40[151]    = ( l_41 [300] & !i[1819]) | ( l_41 [301] &  i[1819]);
assign l_40[152]    = ( l_41 [302] & !i[1819]) | ( l_41 [303] &  i[1819]);
assign l_40[153]    = ( l_41 [304] & !i[1819]) | ( l_41 [305] &  i[1819]);
assign l_40[154]    = ( l_41 [306] & !i[1819]) | ( l_41 [307] &  i[1819]);
assign l_40[155]    = ( l_41 [308] & !i[1819]) | ( l_41 [309] &  i[1819]);
assign l_40[156]    = ( l_41 [310] & !i[1819]) | ( l_41 [311] &  i[1819]);
assign l_40[157]    = ( l_41 [312] & !i[1819]) | ( l_41 [313] &  i[1819]);
assign l_40[158]    = ( l_41 [314] & !i[1819]) | ( l_41 [315] &  i[1819]);
assign l_40[159]    = ( l_41 [316] & !i[1819]) | ( l_41 [317] &  i[1819]);
assign l_40[160]    = ( l_41 [318] & !i[1819]) | ( l_41 [319] &  i[1819]);
assign l_40[161]    = ( l_41 [320] & !i[1819]) | ( l_41 [321] &  i[1819]);
assign l_40[162]    = ( l_41 [322] & !i[1819]) | ( l_41 [323] &  i[1819]);
assign l_40[163]    = ( l_41 [324] & !i[1819]) | ( l_41 [325] &  i[1819]);
assign l_40[164]    = ( l_41 [326] & !i[1819]) | ( l_41 [327] &  i[1819]);
assign l_40[165]    = ( l_41 [328] & !i[1819]) | ( l_41 [329] &  i[1819]);
assign l_40[166]    = ( l_41 [330] & !i[1819]) | ( l_41 [331] &  i[1819]);
assign l_40[167]    = ( l_41 [332] & !i[1819]) | ( l_41 [333] &  i[1819]);
assign l_40[168]    = ( l_41 [334] & !i[1819]) | ( l_41 [335] &  i[1819]);
assign l_40[169]    = ( l_41 [336] & !i[1819]) | ( l_41 [337] &  i[1819]);
assign l_40[170]    = ( l_41 [338] & !i[1819]) | ( l_41 [339] &  i[1819]);
assign l_40[171]    = ( l_41 [340] & !i[1819]) | ( l_41 [341] &  i[1819]);
assign l_40[172]    = ( l_41 [342] & !i[1819]) | ( l_41 [343] &  i[1819]);
assign l_40[173]    = ( l_41 [344] & !i[1819]) | ( l_41 [345] &  i[1819]);
assign l_40[174]    = ( l_41 [346] & !i[1819]) | ( l_41 [347] &  i[1819]);
assign l_40[175]    = ( l_41 [348] & !i[1819]) | ( l_41 [349] &  i[1819]);
assign l_40[176]    = ( l_41 [350] & !i[1819]) | ( l_41 [351] &  i[1819]);
assign l_40[177]    = ( l_41 [352] & !i[1819]) | ( l_41 [353] &  i[1819]);
assign l_40[178]    = ( l_41 [354] & !i[1819]) | ( l_41 [355] &  i[1819]);
assign l_40[179]    = ( l_41 [356] & !i[1819]) | ( l_41 [357] &  i[1819]);
assign l_40[180]    = ( l_41 [358] & !i[1819]) | ( l_41 [359] &  i[1819]);
assign l_40[181]    = ( l_41 [360] & !i[1819]) | ( l_41 [361] &  i[1819]);
assign l_40[182]    = ( l_41 [362] & !i[1819]) | ( l_41 [363] &  i[1819]);
assign l_40[183]    = ( l_41 [364] & !i[1819]) | ( l_41 [365] &  i[1819]);
assign l_40[184]    = ( l_41 [366] & !i[1819]) | ( l_41 [367] &  i[1819]);
assign l_40[185]    = ( l_41 [368] & !i[1819]) | ( l_41 [369] &  i[1819]);
assign l_40[186]    = ( l_41 [370] & !i[1819]) | ( l_41 [371] &  i[1819]);
assign l_40[187]    = ( l_41 [372] & !i[1819]) | ( l_41 [373] &  i[1819]);
assign l_40[188]    = ( l_41 [374] & !i[1819]) | ( l_41 [375] &  i[1819]);
assign l_40[189]    = ( l_41 [376] & !i[1819]) | ( l_41 [377] &  i[1819]);
assign l_40[190]    = ( l_41 [378] & !i[1819]) | ( l_41 [379] &  i[1819]);
assign l_40[191]    = ( l_41 [380] & !i[1819]) | ( l_41 [381] &  i[1819]);
assign l_40[192]    = ( l_41 [382] & !i[1819]) | ( l_41 [383] &  i[1819]);
assign l_40[193]    = ( l_41 [384] & !i[1819]) | ( l_41 [385] &  i[1819]);
assign l_40[194]    = ( l_41 [386] & !i[1819]) | ( l_41 [387] &  i[1819]);
assign l_40[195]    = ( l_41 [388] & !i[1819]) | ( l_41 [389] &  i[1819]);
assign l_40[196]    = ( l_41 [390] & !i[1819]) | ( l_41 [391] &  i[1819]);
assign l_40[197]    = ( l_41 [392] & !i[1819]) | ( l_41 [393] &  i[1819]);
assign l_40[198]    = ( l_41 [394] & !i[1819]) | ( l_41 [395] &  i[1819]);
assign l_40[199]    = ( l_41 [396] & !i[1819]) | ( l_41 [397] &  i[1819]);
assign l_40[200]    = ( l_41 [398] & !i[1819]) | ( l_41 [399] &  i[1819]);
assign l_40[201]    = ( l_41 [400] & !i[1819]) | ( l_41 [401] &  i[1819]);
assign l_40[202]    = ( l_41 [402] & !i[1819]) | ( l_41 [403] &  i[1819]);
assign l_40[203]    = ( l_41 [404] & !i[1819]) | ( l_41 [405] &  i[1819]);
assign l_40[204]    = ( l_41 [406] & !i[1819]) | ( l_41 [407] &  i[1819]);
assign l_40[205]    = ( l_41 [408] & !i[1819]) | ( l_41 [409] &  i[1819]);
assign l_40[206]    = ( l_41 [410] & !i[1819]) | ( l_41 [411] &  i[1819]);
assign l_40[207]    = ( l_41 [412] & !i[1819]) | ( l_41 [413] &  i[1819]);
assign l_40[208]    = ( l_41 [414] & !i[1819]) | ( l_41 [415] &  i[1819]);
assign l_40[209]    = ( l_41 [416] & !i[1819]) | ( l_41 [417] &  i[1819]);
assign l_40[210]    = ( l_41 [418] & !i[1819]) | ( l_41 [419] &  i[1819]);
assign l_40[211]    = ( l_41 [420] & !i[1819]) | ( l_41 [421] &  i[1819]);
assign l_40[212]    = ( l_41 [422] & !i[1819]) | ( l_41 [423] &  i[1819]);
assign l_40[213]    = ( l_41 [424] & !i[1819]) | ( l_41 [425] &  i[1819]);
assign l_40[214]    = ( l_41 [426] & !i[1819]) | ( l_41 [427] &  i[1819]);
assign l_40[215]    = ( l_41 [428] & !i[1819]) | ( l_41 [429] &  i[1819]);
assign l_40[216]    = ( l_41 [430] & !i[1819]) | ( l_41 [431] &  i[1819]);
assign l_40[217]    = ( l_41 [432] & !i[1819]) | ( l_41 [433] &  i[1819]);
assign l_40[218]    = ( l_41 [434] & !i[1819]) | ( l_41 [435] &  i[1819]);
assign l_40[219]    = ( l_41 [436] & !i[1819]) | ( l_41 [437] &  i[1819]);
assign l_40[220]    = ( l_41 [438] & !i[1819]) | ( l_41 [439] &  i[1819]);
assign l_40[221]    = ( l_41 [440] & !i[1819]) | ( l_41 [441] &  i[1819]);
assign l_40[222]    = ( l_41 [442] & !i[1819]) | ( l_41 [443] &  i[1819]);
assign l_40[223]    = ( l_41 [444] & !i[1819]) | ( l_41 [445] &  i[1819]);
assign l_40[224]    = ( l_41 [446] & !i[1819]) | ( l_41 [447] &  i[1819]);
assign l_40[225]    = ( l_41 [448] & !i[1819]) | ( l_41 [449] &  i[1819]);
assign l_40[226]    = ( l_41 [450] & !i[1819]) | ( l_41 [451] &  i[1819]);
assign l_40[227]    = ( l_41 [452] & !i[1819]) | ( l_41 [453] &  i[1819]);
assign l_40[228]    = ( l_41 [454] & !i[1819]) | ( l_41 [455] &  i[1819]);
assign l_40[229]    = ( l_41 [456] & !i[1819]) | ( l_41 [457] &  i[1819]);
assign l_40[230]    = ( l_41 [458] & !i[1819]) | ( l_41 [459] &  i[1819]);
assign l_40[231]    = ( l_41 [460] & !i[1819]) | ( l_41 [461] &  i[1819]);
assign l_40[232]    = ( l_41 [462] & !i[1819]) | ( l_41 [463] &  i[1819]);
assign l_40[233]    = ( l_41 [464] & !i[1819]) | ( l_41 [465] &  i[1819]);
assign l_40[234]    = ( l_41 [466] & !i[1819]) | ( l_41 [467] &  i[1819]);
assign l_40[235]    = ( l_41 [468] & !i[1819]) | ( l_41 [469] &  i[1819]);
assign l_40[236]    = ( l_41 [470] & !i[1819]) | ( l_41 [471] &  i[1819]);
assign l_40[237]    = ( l_41 [472] & !i[1819]) | ( l_41 [473] &  i[1819]);
assign l_40[238]    = ( l_41 [474] & !i[1819]) | ( l_41 [475] &  i[1819]);
assign l_40[239]    = ( l_41 [476] & !i[1819]) | ( l_41 [477] &  i[1819]);
assign l_40[240]    = ( l_41 [478] & !i[1819]) | ( l_41 [479] &  i[1819]);
assign l_40[241]    = ( l_41 [480] & !i[1819]) | ( l_41 [481] &  i[1819]);
assign l_40[242]    = ( l_41 [482] & !i[1819]) | ( l_41 [483] &  i[1819]);
assign l_40[243]    = ( l_41 [484] & !i[1819]) | ( l_41 [485] &  i[1819]);
assign l_40[244]    = ( l_41 [486] & !i[1819]) | ( l_41 [487] &  i[1819]);
assign l_40[245]    = ( l_41 [488] & !i[1819]) | ( l_41 [489] &  i[1819]);
assign l_40[246]    = ( l_41 [490] & !i[1819]) | ( l_41 [491] &  i[1819]);
assign l_40[247]    = ( l_41 [492] & !i[1819]) | ( l_41 [493] &  i[1819]);
assign l_40[248]    = ( l_41 [494] & !i[1819]) | ( l_41 [495] &  i[1819]);
assign l_40[249]    = ( l_41 [496] & !i[1819]) | ( l_41 [497] &  i[1819]);
assign l_40[250]    = ( l_41 [498] & !i[1819]) | ( l_41 [499] &  i[1819]);
assign l_40[251]    = ( l_41 [500] & !i[1819]) | ( l_41 [501] &  i[1819]);
assign l_40[252]    = ( l_41 [502] & !i[1819]) | ( l_41 [503] &  i[1819]);
assign l_40[253]    = ( l_41 [504] & !i[1819]) | ( l_41 [505] &  i[1819]);
assign l_40[254]    = ( l_41 [506] & !i[1819]) | ( l_41 [507] &  i[1819]);
assign l_40[255]    = ( l_41 [508] & !i[1819]) | ( l_41 [509] &  i[1819]);
assign l_40[256]    = ( l_41 [510] & !i[1819]) | ( l_41 [511] &  i[1819]);
assign l_40[257]    = ( l_41 [512] & !i[1819]) | ( l_41 [513] &  i[1819]);
assign l_40[258]    = ( l_41 [514] & !i[1819]) | ( l_41 [515] &  i[1819]);
assign l_40[259]    = ( l_41 [516] & !i[1819]) | ( l_41 [517] &  i[1819]);
assign l_40[260]    = ( l_41 [518] & !i[1819]) | ( l_41 [519] &  i[1819]);
assign l_40[261]    = ( l_41 [520] & !i[1819]) | ( l_41 [521] &  i[1819]);
assign l_40[262]    = ( l_41 [522] & !i[1819]) | ( l_41 [523] &  i[1819]);
assign l_40[263]    = ( l_41 [524] & !i[1819]) | ( l_41 [525] &  i[1819]);
assign l_40[264]    = ( l_41 [526] & !i[1819]) | ( l_41 [527] &  i[1819]);
assign l_40[265]    = ( l_41 [528] & !i[1819]) | ( l_41 [529] &  i[1819]);
assign l_40[266]    = ( l_41 [530] & !i[1819]) | ( l_41 [531] &  i[1819]);
assign l_40[267]    = ( l_41 [532] & !i[1819]) | ( l_41 [533] &  i[1819]);
assign l_40[268]    = ( l_41 [534] & !i[1819]) | ( l_41 [535] &  i[1819]);
assign l_40[269]    = ( l_41 [536] & !i[1819]) | ( l_41 [537] &  i[1819]);
assign l_40[270]    = ( l_41 [538] & !i[1819]) | ( l_41 [539] &  i[1819]);
assign l_40[271]    = ( l_41 [540] & !i[1819]) | ( l_41 [541] &  i[1819]);
assign l_40[272]    = ( l_41 [542] & !i[1819]) | ( l_41 [543] &  i[1819]);
assign l_40[273]    = ( l_41 [544] & !i[1819]) | ( l_41 [545] &  i[1819]);
assign l_40[274]    = ( l_41 [546] & !i[1819]) | ( l_41 [547] &  i[1819]);
assign l_40[275]    = ( l_41 [548] & !i[1819]) | ( l_41 [549] &  i[1819]);
assign l_40[276]    = ( l_41 [550] & !i[1819]) | ( l_41 [551] &  i[1819]);
assign l_40[277]    = ( l_41 [552] & !i[1819]) | ( l_41 [553] &  i[1819]);
assign l_40[278]    = ( l_41 [554] & !i[1819]) | ( l_41 [555] &  i[1819]);
assign l_40[279]    = ( l_41 [556] & !i[1819]) | ( l_41 [557] &  i[1819]);
assign l_40[280]    = ( l_41 [558] & !i[1819]) | ( l_41 [559] &  i[1819]);
assign l_40[281]    = ( l_41 [560] & !i[1819]) | ( l_41 [561] &  i[1819]);
assign l_40[282]    = ( l_41 [562] & !i[1819]) | ( l_41 [563] &  i[1819]);
assign l_40[283]    = ( l_41 [564] & !i[1819]) | ( l_41 [565] &  i[1819]);
assign l_40[284]    = ( l_41 [566] & !i[1819]) | ( l_41 [567] &  i[1819]);
assign l_40[285]    = ( l_41 [568] & !i[1819]) | ( l_41 [569] &  i[1819]);
assign l_40[286]    = ( l_41 [570] & !i[1819]) | ( l_41 [571] &  i[1819]);
assign l_40[287]    = ( l_41 [572] & !i[1819]) | ( l_41 [573] &  i[1819]);
assign l_40[288]    = ( l_41 [574] & !i[1819]) | ( l_41 [575] &  i[1819]);
assign l_40[289]    = ( l_41 [576] & !i[1819]) | ( l_41 [577] &  i[1819]);
assign l_40[290]    = ( l_41 [578] & !i[1819]) | ( l_41 [579] &  i[1819]);
assign l_40[291]    = ( l_41 [580] & !i[1819]) | ( l_41 [581] &  i[1819]);
assign l_40[292]    = ( l_41 [582] & !i[1819]) | ( l_41 [583] &  i[1819]);
assign l_40[293]    = ( l_41 [584] & !i[1819]) | ( l_41 [585] &  i[1819]);
assign l_40[294]    = ( l_41 [586] & !i[1819]) | ( l_41 [587] &  i[1819]);
assign l_40[295]    = ( l_41 [588] & !i[1819]) | ( l_41 [589] &  i[1819]);
assign l_40[296]    = ( l_41 [590] & !i[1819]) | ( l_41 [591] &  i[1819]);
assign l_40[297]    = ( l_41 [592] & !i[1819]) | ( l_41 [593] &  i[1819]);
assign l_40[298]    = ( l_41 [594] & !i[1819]) | ( l_41 [595] &  i[1819]);
assign l_40[299]    = ( l_41 [596] & !i[1819]) | ( l_41 [597] &  i[1819]);
assign l_40[300]    = ( l_41 [598] & !i[1819]) | ( l_41 [599] &  i[1819]);
assign l_40[301]    = ( l_41 [600] & !i[1819]) | ( l_41 [601] &  i[1819]);
assign l_40[302]    = ( l_41 [602] & !i[1819]) | ( l_41 [603] &  i[1819]);
assign l_40[303]    = ( l_41 [604] & !i[1819]) | ( l_41 [605] &  i[1819]);
assign l_40[304]    = ( l_41 [606] & !i[1819]) | ( l_41 [607] &  i[1819]);
assign l_40[305]    = ( l_41 [608] & !i[1819]) | ( l_41 [609] &  i[1819]);
assign l_40[306]    = ( l_41 [610] & !i[1819]) | ( l_41 [611] &  i[1819]);
assign l_40[307]    = ( l_41 [612] & !i[1819]) | ( l_41 [613] &  i[1819]);
assign l_40[308]    = ( l_41 [614] & !i[1819]) | ( l_41 [615] &  i[1819]);
assign l_40[309]    = ( l_41 [616] & !i[1819]) | ( l_41 [617] &  i[1819]);
assign l_40[310]    = ( l_41 [618] & !i[1819]) | ( l_41 [619] &  i[1819]);
assign l_40[311]    = ( l_41 [620] & !i[1819]) | ( l_41 [621] &  i[1819]);
assign l_40[312]    = ( l_41 [622] & !i[1819]) | ( l_41 [623] &  i[1819]);
assign l_40[313]    = ( l_41 [624] & !i[1819]) | ( l_41 [625] &  i[1819]);
assign l_40[314]    = ( l_41 [626] & !i[1819]) | ( l_41 [627] &  i[1819]);
assign l_40[315]    = ( l_41 [628] & !i[1819]) | ( l_41 [629] &  i[1819]);
assign l_40[316]    = ( l_41 [630] & !i[1819]) | ( l_41 [631] &  i[1819]);
assign l_40[317]    = ( l_41 [632] & !i[1819]) | ( l_41 [633] &  i[1819]);
assign l_40[318]    = ( l_41 [634] & !i[1819]) | ( l_41 [635] &  i[1819]);
assign l_40[319]    = ( l_41 [636] & !i[1819]) | ( l_41 [637] &  i[1819]);
assign l_40[320]    = ( l_41 [638] & !i[1819]) | ( l_41 [639] &  i[1819]);
assign l_40[321]    = ( l_41 [640] & !i[1819]) | ( l_41 [641] &  i[1819]);
assign l_40[322]    = ( l_41 [642] & !i[1819]) | ( l_41 [643] &  i[1819]);
assign l_40[323]    = ( l_41 [644] & !i[1819]) | ( l_41 [645] &  i[1819]);
assign l_40[324]    = ( l_41 [646] & !i[1819]) | ( l_41 [647] &  i[1819]);
assign l_40[325]    = ( l_41 [648] & !i[1819]) | ( l_41 [649] &  i[1819]);
assign l_40[326]    = ( l_41 [650] & !i[1819]) | ( l_41 [651] &  i[1819]);
assign l_40[327]    = ( l_41 [652] & !i[1819]) | ( l_41 [653] &  i[1819]);
assign l_40[328]    = ( l_41 [654] & !i[1819]) | ( l_41 [655] &  i[1819]);
assign l_40[329]    = ( l_41 [656] & !i[1819]) | ( l_41 [657] &  i[1819]);
assign l_40[330]    = ( l_41 [658] & !i[1819]) | ( l_41 [659] &  i[1819]);
assign l_40[331]    = ( l_41 [660] & !i[1819]) | ( l_41 [661] &  i[1819]);
assign l_40[332]    = ( l_41 [662] & !i[1819]) | ( l_41 [663] &  i[1819]);
assign l_40[333]    = ( l_41 [664] & !i[1819]) | ( l_41 [665] &  i[1819]);
assign l_40[334]    = ( l_41 [666] & !i[1819]) | ( l_41 [667] &  i[1819]);
assign l_40[335]    = ( l_41 [668] & !i[1819]) | ( l_41 [669] &  i[1819]);
assign l_40[336]    = ( l_41 [670] & !i[1819]) | ( l_41 [671] &  i[1819]);
assign l_40[337]    = ( l_41 [672] & !i[1819]) | ( l_41 [673] &  i[1819]);
assign l_40[338]    = ( l_41 [674] & !i[1819]) | ( l_41 [675] &  i[1819]);
assign l_40[339]    = ( l_41 [676] & !i[1819]) | ( l_41 [677] &  i[1819]);
assign l_40[340]    = ( l_41 [678] & !i[1819]) | ( l_41 [679] &  i[1819]);
assign l_40[341]    = ( l_41 [680] & !i[1819]) | ( l_41 [681] &  i[1819]);
assign l_40[342]    = ( l_41 [682] & !i[1819]) | ( l_41 [683] &  i[1819]);
assign l_40[343]    = ( l_41 [684] & !i[1819]) | ( l_41 [685] &  i[1819]);
assign l_40[344]    = ( l_41 [686] & !i[1819]) | ( l_41 [687] &  i[1819]);
assign l_40[345]    = ( l_41 [688] & !i[1819]) | ( l_41 [689] &  i[1819]);
assign l_40[346]    = ( l_41 [690] & !i[1819]) | ( l_41 [691] &  i[1819]);
assign l_40[347]    = ( l_41 [692] & !i[1819]) | ( l_41 [693] &  i[1819]);
assign l_40[348]    = ( l_41 [694] & !i[1819]) | ( l_41 [695] &  i[1819]);
assign l_40[349]    = ( l_41 [696] & !i[1819]) | ( l_41 [697] &  i[1819]);
assign l_40[350]    = ( l_41 [698] & !i[1819]) | ( l_41 [699] &  i[1819]);
assign l_40[351]    = ( l_41 [700] & !i[1819]) | ( l_41 [701] &  i[1819]);
assign l_40[352]    = ( l_41 [702] & !i[1819]) | ( l_41 [703] &  i[1819]);
assign l_40[353]    = ( l_41 [704] & !i[1819]) | ( l_41 [705] &  i[1819]);
assign l_40[354]    = ( l_41 [706] & !i[1819]) | ( l_41 [707] &  i[1819]);
assign l_40[355]    = ( l_41 [708] & !i[1819]) | ( l_41 [709] &  i[1819]);
assign l_40[356]    = ( l_41 [710] & !i[1819]) | ( l_41 [711] &  i[1819]);
assign l_40[357]    = ( l_41 [712] & !i[1819]) | ( l_41 [713] &  i[1819]);
assign l_40[358]    = ( l_41 [714] & !i[1819]) | ( l_41 [715] &  i[1819]);
assign l_40[359]    = ( l_41 [716] & !i[1819]) | ( l_41 [717] &  i[1819]);
assign l_40[360]    = ( l_41 [718] & !i[1819]) | ( l_41 [719] &  i[1819]);
assign l_40[361]    = ( l_41 [720] & !i[1819]) | ( l_41 [721] &  i[1819]);
assign l_40[362]    = ( l_41 [722] & !i[1819]) | ( l_41 [723] &  i[1819]);
assign l_40[363]    = ( l_41 [724] & !i[1819]) | ( l_41 [725] &  i[1819]);
assign l_40[364]    = ( l_41 [726] & !i[1819]) | ( l_41 [727] &  i[1819]);
assign l_40[365]    = ( l_41 [728] & !i[1819]) | ( l_41 [729] &  i[1819]);
assign l_40[366]    = ( l_41 [730] & !i[1819]) | ( l_41 [731] &  i[1819]);
assign l_40[367]    = ( l_41 [732] & !i[1819]) | ( l_41 [733] &  i[1819]);
assign l_40[368]    = ( l_41 [734] & !i[1819]) | ( l_41 [735] &  i[1819]);
assign l_40[369]    = ( l_41 [736] & !i[1819]) | ( l_41 [737] &  i[1819]);
assign l_40[370]    = ( l_41 [738] & !i[1819]) | ( l_41 [739] &  i[1819]);
assign l_40[371]    = ( l_41 [740] & !i[1819]) | ( l_41 [741] &  i[1819]);
assign l_40[372]    = ( l_41 [742] & !i[1819]) | ( l_41 [743] &  i[1819]);
assign l_40[373]    = ( l_41 [744] & !i[1819]) | ( l_41 [745] &  i[1819]);
assign l_40[374]    = ( l_41 [746] & !i[1819]) | ( l_41 [747] &  i[1819]);
assign l_40[375]    = ( l_41 [748] & !i[1819]) | ( l_41 [749] &  i[1819]);
assign l_40[376]    = ( l_41 [750] & !i[1819]) | ( l_41 [751] &  i[1819]);
assign l_40[377]    = ( l_41 [752] & !i[1819]) | ( l_41 [753] &  i[1819]);
assign l_40[378]    = ( l_41 [754] & !i[1819]) | ( l_41 [755] &  i[1819]);
assign l_40[379]    = ( l_41 [756] & !i[1819]) | ( l_41 [757] &  i[1819]);
assign l_40[380]    = ( l_41 [758] & !i[1819]) | ( l_41 [759] &  i[1819]);
assign l_40[381]    = ( l_41 [760] & !i[1819]) | ( l_41 [761] &  i[1819]);
assign l_40[382]    = ( l_41 [762] & !i[1819]) | ( l_41 [763] &  i[1819]);
assign l_40[383]    = ( l_41 [764] & !i[1819]) | ( l_41 [765] &  i[1819]);
assign l_40[384]    = ( l_41 [766] & !i[1819]) | ( l_41 [767] &  i[1819]);
assign l_40[385]    = ( l_41 [768] & !i[1819]) | ( l_41 [769] &  i[1819]);
assign l_40[386]    = ( l_41 [770] & !i[1819]) | ( l_41 [771] &  i[1819]);
assign l_40[387]    = ( l_41 [772] & !i[1819]) | ( l_41 [773] &  i[1819]);
assign l_40[388]    = ( l_41 [774] & !i[1819]) | ( l_41 [775] &  i[1819]);
assign l_40[389]    = ( l_41 [776] & !i[1819]) | ( l_41 [777] &  i[1819]);
assign l_40[390]    = ( l_41 [778] & !i[1819]) | ( l_41 [779] &  i[1819]);
assign l_40[391]    = ( l_41 [780] & !i[1819]) | ( l_41 [781] &  i[1819]);
assign l_40[392]    = ( l_41 [782] & !i[1819]) | ( l_41 [783] &  i[1819]);
assign l_40[393]    = ( l_41 [784] & !i[1819]) | ( l_41 [785] &  i[1819]);
assign l_40[394]    = ( l_41 [786] & !i[1819]) | ( l_41 [787] &  i[1819]);
assign l_40[395]    = ( l_41 [788] & !i[1819]) | ( l_41 [789] &  i[1819]);
assign l_40[396]    = ( l_41 [790] & !i[1819]) | ( l_41 [791] &  i[1819]);
assign l_40[397]    = ( l_41 [792] & !i[1819]) | ( l_41 [793] &  i[1819]);
assign l_40[398]    = ( l_41 [794] & !i[1819]) | ( l_41 [795] &  i[1819]);
assign l_40[399]    = ( l_41 [796] & !i[1819]) | ( l_41 [797] &  i[1819]);
assign l_40[400]    = ( l_41 [798] & !i[1819]) | ( l_41 [799] &  i[1819]);
assign l_40[401]    = ( l_41 [800] & !i[1819]) | ( l_41 [801] &  i[1819]);
assign l_40[402]    = ( l_41 [802] & !i[1819]) | ( l_41 [803] &  i[1819]);
assign l_40[403]    = ( l_41 [804] & !i[1819]) | ( l_41 [805] &  i[1819]);
assign l_40[404]    = ( l_41 [806] & !i[1819]) | ( l_41 [807] &  i[1819]);
assign l_40[405]    = ( l_41 [808] & !i[1819]) | ( l_41 [809] &  i[1819]);
assign l_40[406]    = ( l_41 [810] & !i[1819]) | ( l_41 [811] &  i[1819]);
assign l_40[407]    = ( l_41 [812] & !i[1819]) | ( l_41 [813] &  i[1819]);
assign l_40[408]    = ( l_41 [814] & !i[1819]) | ( l_41 [815] &  i[1819]);
assign l_40[409]    = ( l_41 [816] & !i[1819]) | ( l_41 [817] &  i[1819]);
assign l_40[410]    = ( l_41 [818] & !i[1819]) | ( l_41 [819] &  i[1819]);
assign l_40[411]    = ( l_41 [820] & !i[1819]) | ( l_41 [821] &  i[1819]);
assign l_40[412]    = ( l_41 [822] & !i[1819]) | ( l_41 [823] &  i[1819]);
assign l_40[413]    = ( l_41 [824] & !i[1819]) | ( l_41 [825] &  i[1819]);
assign l_40[414]    = ( l_41 [826] & !i[1819]) | ( l_41 [827] &  i[1819]);
assign l_40[415]    = ( l_41 [828] & !i[1819]) | ( l_41 [829] &  i[1819]);
assign l_40[416]    = ( l_41 [830] & !i[1819]) | ( l_41 [831] &  i[1819]);
assign l_40[417]    = ( l_41 [832] & !i[1819]) | ( l_41 [833] &  i[1819]);
assign l_40[418]    = ( l_41 [834] & !i[1819]) | ( l_41 [835] &  i[1819]);
assign l_40[419]    = ( l_41 [836] & !i[1819]) | ( l_41 [837] &  i[1819]);
assign l_40[420]    = ( l_41 [838] & !i[1819]) | ( l_41 [839] &  i[1819]);
assign l_40[421]    = ( l_41 [840] & !i[1819]) | ( l_41 [841] &  i[1819]);
assign l_40[422]    = ( l_41 [842] & !i[1819]) | ( l_41 [843] &  i[1819]);
assign l_40[423]    = ( l_41 [844] & !i[1819]) | ( l_41 [845] &  i[1819]);
assign l_40[424]    = ( l_41 [846] & !i[1819]) | ( l_41 [847] &  i[1819]);
assign l_40[425]    = ( l_41 [848] & !i[1819]) | ( l_41 [849] &  i[1819]);
assign l_40[426]    = ( l_41 [850] & !i[1819]) | ( l_41 [851] &  i[1819]);
assign l_40[427]    = ( l_41 [852] & !i[1819]) | ( l_41 [853] &  i[1819]);
assign l_40[428]    = ( l_41 [854] & !i[1819]) | ( l_41 [855] &  i[1819]);
assign l_40[429]    = ( l_41 [856] & !i[1819]) | ( l_41 [857] &  i[1819]);
assign l_40[430]    = ( l_41 [858] & !i[1819]) | ( l_41 [859] &  i[1819]);
assign l_40[431]    = ( l_41 [860] & !i[1819]) | ( l_41 [861] &  i[1819]);
assign l_40[432]    = ( l_41 [862] & !i[1819]) | ( l_41 [863] &  i[1819]);
assign l_40[433]    = ( l_41 [864] & !i[1819]) | ( l_41 [865] &  i[1819]);
assign l_40[434]    = ( l_41 [866] & !i[1819]) | ( l_41 [867] &  i[1819]);
assign l_40[435]    = ( l_41 [868] & !i[1819]) | ( l_41 [869] &  i[1819]);
assign l_40[436]    = ( l_41 [870] & !i[1819]) | ( l_41 [871] &  i[1819]);
assign l_40[437]    = ( l_41 [872] & !i[1819]) | ( l_41 [873] &  i[1819]);
assign l_40[438]    = ( l_41 [874] & !i[1819]) | ( l_41 [875] &  i[1819]);
assign l_40[439]    = ( l_41 [876] & !i[1819]) | ( l_41 [877] &  i[1819]);
assign l_40[440]    = ( l_41 [878] & !i[1819]) | ( l_41 [879] &  i[1819]);
assign l_40[441]    = ( l_41 [880] & !i[1819]) | ( l_41 [881] &  i[1819]);
assign l_40[442]    = ( l_41 [882] & !i[1819]) | ( l_41 [883] &  i[1819]);
assign l_40[443]    = ( l_41 [884] & !i[1819]) | ( l_41 [885] &  i[1819]);
assign l_40[444]    = ( l_41 [886] & !i[1819]) | ( l_41 [887] &  i[1819]);
assign l_40[445]    = ( l_41 [888] & !i[1819]) | ( l_41 [889] &  i[1819]);
assign l_40[446]    = ( l_41 [890] & !i[1819]) | ( l_41 [891] &  i[1819]);
assign l_40[447]    = ( l_41 [892] & !i[1819]) | ( l_41 [893] &  i[1819]);
assign l_40[448]    = ( l_41 [894] & !i[1819]) | ( l_41 [895] &  i[1819]);
assign l_40[449]    = ( l_41 [896] & !i[1819]) | ( l_41 [897] &  i[1819]);
assign l_40[450]    = ( l_41 [898] & !i[1819]) | ( l_41 [899] &  i[1819]);
assign l_40[451]    = ( l_41 [900] & !i[1819]) | ( l_41 [901] &  i[1819]);
assign l_40[452]    = ( l_41 [902] & !i[1819]) | ( l_41 [903] &  i[1819]);
assign l_40[453]    = ( l_41 [904] & !i[1819]) | ( l_41 [905] &  i[1819]);
assign l_40[454]    = ( l_41 [906] & !i[1819]) | ( l_41 [907] &  i[1819]);
assign l_40[455]    = ( l_41 [908] & !i[1819]) | ( l_41 [909] &  i[1819]);
assign l_40[456]    = ( l_41 [910] & !i[1819]) | ( l_41 [911] &  i[1819]);
assign l_40[457]    = ( l_41 [912] & !i[1819]) | ( l_41 [913] &  i[1819]);
assign l_40[458]    = ( l_41 [914] & !i[1819]) | ( l_41 [915] &  i[1819]);
assign l_40[459]    = ( l_41 [916] & !i[1819]) | ( l_41 [917] &  i[1819]);
assign l_40[460]    = ( l_41 [918] & !i[1819]) | ( l_41 [919] &  i[1819]);
assign l_40[461]    = ( l_41 [920] & !i[1819]) | ( l_41 [921] &  i[1819]);
assign l_40[462]    = ( l_41 [922] & !i[1819]) | ( l_41 [923] &  i[1819]);
assign l_40[463]    = ( l_41 [924] & !i[1819]) | ( l_41 [925] &  i[1819]);
assign l_40[464]    = ( l_41 [926] & !i[1819]) | ( l_41 [927] &  i[1819]);
assign l_40[465]    = ( l_41 [928] & !i[1819]) | ( l_41 [929] &  i[1819]);
assign l_40[466]    = ( l_41 [930] & !i[1819]) | ( l_41 [931] &  i[1819]);
assign l_40[467]    = ( l_41 [932] & !i[1819]) | ( l_41 [933] &  i[1819]);
assign l_40[468]    = ( l_41 [934] & !i[1819]) | ( l_41 [935] &  i[1819]);
assign l_40[469]    = ( l_41 [936] & !i[1819]) | ( l_41 [937] &  i[1819]);
assign l_40[470]    = ( l_41 [938] & !i[1819]) | ( l_41 [939] &  i[1819]);
assign l_40[471]    = ( l_41 [940] & !i[1819]) | ( l_41 [941] &  i[1819]);
assign l_40[472]    = ( l_41 [942] & !i[1819]) | ( l_41 [943] &  i[1819]);
assign l_40[473]    = ( l_41 [944] & !i[1819]) | ( l_41 [945] &  i[1819]);
assign l_40[474]    = ( l_41 [946] & !i[1819]) | ( l_41 [947] &  i[1819]);
assign l_40[475]    = ( l_41 [948] & !i[1819]) | ( l_41 [949] &  i[1819]);
assign l_40[476]    = ( l_41 [950] & !i[1819]) | ( l_41 [951] &  i[1819]);
assign l_40[477]    = ( l_41 [952] & !i[1819]) | ( l_41 [953] &  i[1819]);
assign l_40[478]    = ( l_41 [954] & !i[1819]) | ( l_41 [955] &  i[1819]);
assign l_40[479]    = ( l_41 [956] & !i[1819]) | ( l_41 [957] &  i[1819]);
assign l_40[480]    = ( l_41 [958] & !i[1819]) | ( l_41 [959] &  i[1819]);
assign l_40[481]    = ( l_41 [960] & !i[1819]) | ( l_41 [961] &  i[1819]);
assign l_40[482]    = ( l_41 [962] & !i[1819]) | ( l_41 [963] &  i[1819]);
assign l_40[483]    = ( l_41 [964] & !i[1819]) | ( l_41 [965] &  i[1819]);
assign l_40[484]    = ( l_41 [966] & !i[1819]) | ( l_41 [967] &  i[1819]);
assign l_40[485]    = ( l_41 [968] & !i[1819]) | ( l_41 [969] &  i[1819]);
assign l_40[486]    = ( l_41 [970] & !i[1819]) | ( l_41 [971] &  i[1819]);
assign l_40[487]    = ( l_41 [972] & !i[1819]) | ( l_41 [973] &  i[1819]);
assign l_40[488]    = ( l_41 [974] & !i[1819]) | ( l_41 [975] &  i[1819]);
assign l_40[489]    = ( l_41 [976] & !i[1819]) | ( l_41 [977] &  i[1819]);
assign l_40[490]    = ( l_41 [978] & !i[1819]) | ( l_41 [979] &  i[1819]);
assign l_40[491]    = ( l_41 [980] & !i[1819]) | ( l_41 [981] &  i[1819]);
assign l_40[492]    = ( l_41 [982] & !i[1819]) | ( l_41 [983] &  i[1819]);
assign l_40[493]    = ( l_41 [984] & !i[1819]) | ( l_41 [985] &  i[1819]);
assign l_40[494]    = ( l_41 [986] & !i[1819]) | ( l_41 [987] &  i[1819]);
assign l_40[495]    = ( l_41 [988] & !i[1819]) | ( l_41 [989] &  i[1819]);
assign l_40[496]    = ( l_41 [990] & !i[1819]) | ( l_41 [991] &  i[1819]);
assign l_40[497]    = ( l_41 [992] & !i[1819]) | ( l_41 [993] &  i[1819]);
assign l_40[498]    = ( l_41 [994] & !i[1819]) | ( l_41 [995] &  i[1819]);
assign l_40[499]    = ( l_41 [996] & !i[1819]) | ( l_41 [997] &  i[1819]);
assign l_40[500]    = ( l_41 [998] & !i[1819]) | ( l_41 [999] &  i[1819]);
assign l_40[501]    = ( l_41 [1000] & !i[1819]) | ( l_41 [1001] &  i[1819]);
assign l_40[502]    = ( l_41 [1002] & !i[1819]) | ( l_41 [1003] &  i[1819]);
assign l_40[503]    = ( l_41 [1004] & !i[1819]) | ( l_41 [1005] &  i[1819]);
assign l_40[504]    = ( l_41 [1006] & !i[1819]) | ( l_41 [1007] &  i[1819]);
assign l_40[505]    = ( l_41 [1008] & !i[1819]) | ( l_41 [1009] &  i[1819]);
assign l_40[506]    = ( l_41 [1010] & !i[1819]) | ( l_41 [1011] &  i[1819]);
assign l_40[507]    = ( l_41 [1012] & !i[1819]) | ( l_41 [1013] &  i[1819]);
assign l_40[508]    = ( l_41 [1014] & !i[1819]) | ( l_41 [1015] &  i[1819]);
assign l_40[509]    = ( l_41 [1016] & !i[1819]) | ( l_41 [1017] &  i[1819]);
assign l_40[510]    = ( l_41 [1018] & !i[1819]) | ( l_41 [1019] &  i[1819]);
assign l_40[511]    = ( l_41 [1020] & !i[1819]) | ( l_41 [1021] &  i[1819]);
assign l_40[512]    = ( l_41 [1022] & !i[1819]) | ( l_41 [1023] &  i[1819]);
assign l_40[513]    = ( l_41 [1024] & !i[1819]) | ( l_41 [1025] &  i[1819]);
assign l_40[514]    = ( l_41 [1026] & !i[1819]) | ( l_41 [1027] &  i[1819]);
assign l_40[515]    = ( l_41 [1028] & !i[1819]) | ( l_41 [1029] &  i[1819]);
assign l_40[516]    = ( l_41 [1030] & !i[1819]) | ( l_41 [1031] &  i[1819]);
assign l_40[517]    = ( l_41 [1032] & !i[1819]) | ( l_41 [1033] &  i[1819]);
assign l_40[518]    = ( l_41 [1034] & !i[1819]) | ( l_41 [1035] &  i[1819]);
assign l_40[519]    = ( l_41 [1036] & !i[1819]) | ( l_41 [1037] &  i[1819]);
assign l_40[520]    = ( l_41 [1038] & !i[1819]) | ( l_41 [1039] &  i[1819]);
assign l_40[521]    = ( l_41 [1040] & !i[1819]) | ( l_41 [1041] &  i[1819]);
assign l_40[522]    = ( l_41 [1042] & !i[1819]) | ( l_41 [1043] &  i[1819]);
assign l_40[523]    = ( l_41 [1044] & !i[1819]) | ( l_41 [1045] &  i[1819]);
assign l_40[524]    = ( l_41 [1046] & !i[1819]) | ( l_41 [1047] &  i[1819]);
assign l_40[525]    = ( l_41 [1048] & !i[1819]) | ( l_41 [1049] &  i[1819]);
assign l_40[526]    = ( l_41 [1050] & !i[1819]) | ( l_41 [1051] &  i[1819]);
assign l_40[527]    = ( l_41 [1052] & !i[1819]) | ( l_41 [1053] &  i[1819]);
assign l_40[528]    = ( l_41 [1054] & !i[1819]) | ( l_41 [1055] &  i[1819]);
assign l_40[529]    = ( l_41 [1056] & !i[1819]) | ( l_41 [1057] &  i[1819]);
assign l_40[530]    = ( l_41 [1058] & !i[1819]) | ( l_41 [1059] &  i[1819]);
assign l_40[531]    = ( l_41 [1060] & !i[1819]) | ( l_41 [1061] &  i[1819]);
assign l_40[532]    = ( l_41 [1062] & !i[1819]) | ( l_41 [1063] &  i[1819]);
assign l_40[533]    = ( l_41 [1064] & !i[1819]) | ( l_41 [1065] &  i[1819]);
assign l_40[534]    = ( l_41 [1066] & !i[1819]) | ( l_41 [1067] &  i[1819]);
assign l_40[535]    = ( l_41 [1068] & !i[1819]) | ( l_41 [1069] &  i[1819]);
assign l_40[536]    = ( l_41 [1070] & !i[1819]) | ( l_41 [1071] &  i[1819]);
assign l_40[537]    = ( l_41 [1072] & !i[1819]) | ( l_41 [1073] &  i[1819]);
assign l_40[538]    = ( l_41 [1074] & !i[1819]) | ( l_41 [1075] &  i[1819]);
assign l_40[539]    = ( l_41 [1076] & !i[1819]) | ( l_41 [1077] &  i[1819]);
assign l_40[540]    = ( l_41 [1078] & !i[1819]) | ( l_41 [1079] &  i[1819]);
assign l_40[541]    = ( l_41 [1080] & !i[1819]) | ( l_41 [1081] &  i[1819]);
assign l_40[542]    = ( l_41 [1082] & !i[1819]) | ( l_41 [1083] &  i[1819]);
assign l_40[543]    = ( l_41 [1084] & !i[1819]) | ( l_41 [1085] &  i[1819]);
assign l_40[544]    = ( l_41 [1086] & !i[1819]) | ( l_41 [1087] &  i[1819]);
assign l_40[545]    = ( l_41 [1088] & !i[1819]) | ( l_41 [1089] &  i[1819]);
assign l_40[546]    = ( l_41 [1090] & !i[1819]) | ( l_41 [1091] &  i[1819]);
assign l_40[547]    = ( l_41 [1092] & !i[1819]) | ( l_41 [1093] &  i[1819]);
assign l_40[548]    = ( l_41 [1094] & !i[1819]) | ( l_41 [1095] &  i[1819]);
assign l_40[549]    = ( l_41 [1096] & !i[1819]) | ( l_41 [1097] &  i[1819]);
assign l_40[550]    = ( l_41 [1098] & !i[1819]) | ( l_41 [1099] &  i[1819]);
assign l_40[551]    = ( l_41 [1100] & !i[1819]) | ( l_41 [1101] &  i[1819]);
assign l_40[552]    = ( l_41 [1102] & !i[1819]) | ( l_41 [1103] &  i[1819]);
assign l_40[553]    = ( l_41 [1104] & !i[1819]) | ( l_41 [1105] &  i[1819]);
assign l_40[554]    = ( l_41 [1106] & !i[1819]) | ( l_41 [1107] &  i[1819]);
assign l_40[555]    = ( l_41 [1108] & !i[1819]) | ( l_41 [1109] &  i[1819]);
assign l_40[556]    = ( l_41 [1110] & !i[1819]) | ( l_41 [1111] &  i[1819]);
assign l_40[557]    = ( l_41 [1112] & !i[1819]) | ( l_41 [1113] &  i[1819]);
assign l_40[558]    = ( l_41 [1114] & !i[1819]) | ( l_41 [1115] &  i[1819]);
assign l_40[559]    = ( l_41 [1116] & !i[1819]) | ( l_41 [1117] &  i[1819]);
assign l_40[560]    = ( l_41 [1118] & !i[1819]) | ( l_41 [1119] &  i[1819]);
assign l_40[561]    = ( l_41 [1120] & !i[1819]) | ( l_41 [1121] &  i[1819]);
assign l_40[562]    = ( l_41 [1122] & !i[1819]) | ( l_41 [1123] &  i[1819]);
assign l_40[563]    = ( l_41 [1124] & !i[1819]) | ( l_41 [1125] &  i[1819]);
assign l_40[564]    = ( l_41 [1126] & !i[1819]) | ( l_41 [1127] &  i[1819]);
assign l_40[565]    = ( l_41 [1128] & !i[1819]) | ( l_41 [1129] &  i[1819]);
assign l_40[566]    = ( l_41 [1130] & !i[1819]) | ( l_41 [1131] &  i[1819]);
assign l_40[567]    = ( l_41 [1132] & !i[1819]) | ( l_41 [1133] &  i[1819]);
assign l_40[568]    = ( l_41 [1134] & !i[1819]) | ( l_41 [1135] &  i[1819]);
assign l_40[569]    = ( l_41 [1136] & !i[1819]) | ( l_41 [1137] &  i[1819]);
assign l_40[570]    = ( l_41 [1138] & !i[1819]) | ( l_41 [1139] &  i[1819]);
assign l_40[571]    = ( l_41 [1140] & !i[1819]) | ( l_41 [1141] &  i[1819]);
assign l_40[572]    = ( l_41 [1142] & !i[1819]) | ( l_41 [1143] &  i[1819]);
assign l_40[573]    = ( l_41 [1144] & !i[1819]) | ( l_41 [1145] &  i[1819]);
assign l_40[574]    = ( l_41 [1146] & !i[1819]) | ( l_41 [1147] &  i[1819]);
assign l_40[575]    = ( l_41 [1148] & !i[1819]) | ( l_41 [1149] &  i[1819]);
assign l_40[576]    = ( l_41 [1150] & !i[1819]) | ( l_41 [1151] &  i[1819]);
assign l_40[577]    = ( l_41 [1152] & !i[1819]) | ( l_41 [1153] &  i[1819]);
assign l_40[578]    = ( l_41 [1154] & !i[1819]) | ( l_41 [1155] &  i[1819]);
assign l_40[579]    = ( l_41 [1156] & !i[1819]) | ( l_41 [1157] &  i[1819]);
assign l_40[580]    = ( l_41 [1158] & !i[1819]) | ( l_41 [1159] &  i[1819]);
assign l_40[581]    = ( l_41 [1160] & !i[1819]) | ( l_41 [1161] &  i[1819]);
assign l_40[582]    = ( l_41 [1162] & !i[1819]) | ( l_41 [1163] &  i[1819]);
assign l_40[583]    = ( l_41 [1164] & !i[1819]) | ( l_41 [1165] &  i[1819]);
assign l_40[584]    = ( l_41 [1166] & !i[1819]) | ( l_41 [1167] &  i[1819]);
assign l_40[585]    = ( l_41 [1168] & !i[1819]) | ( l_41 [1169] &  i[1819]);
assign l_40[586]    = ( l_41 [1170] & !i[1819]) | ( l_41 [1171] &  i[1819]);
assign l_40[587]    = ( l_41 [1172] & !i[1819]) | ( l_41 [1173] &  i[1819]);
assign l_40[588]    = ( l_41 [1174] & !i[1819]) | ( l_41 [1175] &  i[1819]);
assign l_40[589]    = ( l_41 [1176] & !i[1819]) | ( l_41 [1177] &  i[1819]);
assign l_40[590]    = ( l_41 [1178] & !i[1819]) | ( l_41 [1179] &  i[1819]);
assign l_40[591]    = ( l_41 [1180] & !i[1819]) | ( l_41 [1181] &  i[1819]);
assign l_40[592]    = ( l_41 [1182] & !i[1819]) | ( l_41 [1183] &  i[1819]);
assign l_40[593]    = ( l_41 [1184] & !i[1819]) | ( l_41 [1185] &  i[1819]);
assign l_40[594]    = ( l_41 [1186] & !i[1819]) | ( l_41 [1187] &  i[1819]);
assign l_40[595]    = ( l_41 [1188] & !i[1819]) | ( l_41 [1189] &  i[1819]);
assign l_40[596]    = ( l_41 [1190] & !i[1819]) | ( l_41 [1191] &  i[1819]);
assign l_40[597]    = ( l_41 [1192] & !i[1819]) | ( l_41 [1193] &  i[1819]);
assign l_40[598]    = ( l_41 [1194] & !i[1819]) | ( l_41 [1195] &  i[1819]);
assign l_40[599]    = ( l_41 [1196] & !i[1819]) | ( l_41 [1197] &  i[1819]);
assign l_40[600]    = ( l_41 [1198] & !i[1819]) | ( l_41 [1199] &  i[1819]);
assign l_40[601]    = ( l_41 [1200] & !i[1819]) | ( l_41 [1201] &  i[1819]);
assign l_40[602]    = ( l_41 [1202] & !i[1819]) | ( l_41 [1203] &  i[1819]);
assign l_40[603]    = ( l_41 [1204] & !i[1819]) | ( l_41 [1205] &  i[1819]);
assign l_40[604]    = ( l_41 [1206] & !i[1819]) | ( l_41 [1207] &  i[1819]);
assign l_40[605]    = ( l_41 [1208] & !i[1819]) | ( l_41 [1209] &  i[1819]);
assign l_40[606]    = ( l_41 [1210] & !i[1819]) | ( l_41 [1211] &  i[1819]);
assign l_40[607]    = ( l_41 [1212] & !i[1819]) | ( l_41 [1213] &  i[1819]);
assign l_40[608]    = ( l_41 [1214] & !i[1819]) | ( l_41 [1215] &  i[1819]);
assign l_40[609]    = ( l_41 [1216] & !i[1819]) | ( l_41 [1217] &  i[1819]);
assign l_40[610]    = ( l_41 [1218] & !i[1819]) | ( l_41 [1219] &  i[1819]);
assign l_40[611]    = ( l_41 [1220] & !i[1819]) | ( l_41 [1221] &  i[1819]);
assign l_40[612]    = ( l_41 [1222] & !i[1819]) | ( l_41 [1223] &  i[1819]);
assign l_40[613]    = ( l_41 [1224] & !i[1819]) | ( l_41 [1225] &  i[1819]);
assign l_40[614]    = ( l_41 [1226] & !i[1819]) | ( l_41 [1227] &  i[1819]);
assign l_40[615]    = ( l_41 [1228] & !i[1819]) | ( l_41 [1229] &  i[1819]);
assign l_40[616]    = ( l_41 [1230] & !i[1819]) | ( l_41 [1231] &  i[1819]);
assign l_40[617]    = ( l_41 [1232] & !i[1819]) | ( l_41 [1233] &  i[1819]);
assign l_40[618]    = ( l_41 [1234] & !i[1819]) | ( l_41 [1235] &  i[1819]);
assign l_40[619]    = ( l_41 [1236] & !i[1819]) | ( l_41 [1237] &  i[1819]);
assign l_40[620]    = ( l_41 [1238] & !i[1819]) | ( l_41 [1239] &  i[1819]);
assign l_40[621]    = ( l_41 [1240] & !i[1819]) | ( l_41 [1241] &  i[1819]);
assign l_40[622]    = ( l_41 [1242] & !i[1819]) | ( l_41 [1243] &  i[1819]);
assign l_40[623]    = ( l_41 [1244] & !i[1819]) | ( l_41 [1245] &  i[1819]);
assign l_40[624]    = ( l_41 [1246] & !i[1819]) | ( l_41 [1247] &  i[1819]);
assign l_40[625]    = ( l_41 [1248] & !i[1819]) | ( l_41 [1249] &  i[1819]);
assign l_40[626]    = ( l_41 [1250] & !i[1819]) | ( l_41 [1251] &  i[1819]);
assign l_40[627]    = ( l_41 [1252] & !i[1819]) | ( l_41 [1253] &  i[1819]);
assign l_40[628]    = ( l_41 [1254] & !i[1819]) | ( l_41 [1255] &  i[1819]);
assign l_40[629]    = ( l_41 [1256] & !i[1819]) | ( l_41 [1257] &  i[1819]);
assign l_40[630]    = ( l_41 [1258] & !i[1819]) | ( l_41 [1259] &  i[1819]);
assign l_40[631]    = ( l_41 [1260] & !i[1819]) | ( l_41 [1261] &  i[1819]);
assign l_40[632]    = ( l_41 [1262] & !i[1819]) | ( l_41 [1263] &  i[1819]);
assign l_40[633]    = ( l_41 [1264] & !i[1819]) | ( l_41 [1265] &  i[1819]);
assign l_40[634]    = ( l_41 [1266] & !i[1819]) | ( l_41 [1267] &  i[1819]);
assign l_40[635]    = ( l_41 [1268] & !i[1819]) | ( l_41 [1269] &  i[1819]);
assign l_40[636]    = ( l_41 [1270] & !i[1819]) | ( l_41 [1271] &  i[1819]);
assign l_40[637]    = ( l_41 [1272] & !i[1819]) | ( l_41 [1273] &  i[1819]);
assign l_40[638]    = ( l_41 [1274] & !i[1819]) | ( l_41 [1275] &  i[1819]);
assign l_40[639]    = ( l_41 [1276] & !i[1819]) | ( l_41 [1277] &  i[1819]);
assign l_40[640]    = ( l_41 [1278] & !i[1819]) | ( l_41 [1279] &  i[1819]);
assign l_40[641]    = ( l_41 [1280] & !i[1819]) | ( l_41 [1281] &  i[1819]);
assign l_40[642]    = ( l_41 [1282] & !i[1819]) | ( l_41 [1283] &  i[1819]);
assign l_40[643]    = ( l_41 [1284] & !i[1819]) | ( l_41 [1285] &  i[1819]);
assign l_40[644]    = ( l_41 [1286] & !i[1819]) | ( l_41 [1287] &  i[1819]);
assign l_40[645]    = ( l_41 [1288] & !i[1819]) | ( l_41 [1289] &  i[1819]);
assign l_40[646]    = ( l_41 [1290] & !i[1819]) | ( l_41 [1291] &  i[1819]);
assign l_40[647]    = ( l_41 [1292] & !i[1819]) | ( l_41 [1293] &  i[1819]);
assign l_40[648]    = ( l_41 [1294] & !i[1819]) | ( l_41 [1295] &  i[1819]);
assign l_40[649]    = ( l_41 [1296] & !i[1819]) | ( l_41 [1297] &  i[1819]);
assign l_40[650]    = ( l_41 [1298] & !i[1819]) | ( l_41 [1299] &  i[1819]);
assign l_40[651]    = ( l_41 [1300] & !i[1819]) | ( l_41 [1301] &  i[1819]);
assign l_40[652]    = ( l_41 [1302] & !i[1819]) | ( l_41 [1303] &  i[1819]);
assign l_40[653]    = ( l_41 [1304] & !i[1819]) | ( l_41 [1305] &  i[1819]);
assign l_40[654]    = ( l_41 [1306] & !i[1819]) | ( l_41 [1307] &  i[1819]);
assign l_40[655]    = ( l_41 [1308] & !i[1819]) | ( l_41 [1309] &  i[1819]);
assign l_40[656]    = ( l_41 [1310] & !i[1819]) | ( l_41 [1311] &  i[1819]);
assign l_40[657]    = ( l_41 [1312] & !i[1819]) | ( l_41 [1313] &  i[1819]);
assign l_40[658]    = ( l_41 [1314] & !i[1819]) | ( l_41 [1315] &  i[1819]);
assign l_40[659]    = ( l_41 [1316] & !i[1819]) | ( l_41 [1317] &  i[1819]);
assign l_40[660]    = ( l_41 [1318] & !i[1819]) | ( l_41 [1319] &  i[1819]);
assign l_40[661]    = ( l_41 [1320] & !i[1819]) | ( l_41 [1321] &  i[1819]);
assign l_40[662]    = ( l_41 [1322] & !i[1819]) | ( l_41 [1323] &  i[1819]);
assign l_40[663]    = ( l_41 [1324] & !i[1819]) | ( l_41 [1325] &  i[1819]);
assign l_40[664]    = ( l_41 [1326] & !i[1819]) | ( l_41 [1327] &  i[1819]);
assign l_40[665]    = ( l_41 [1328] & !i[1819]) | ( l_41 [1329] &  i[1819]);
assign l_40[666]    = ( l_41 [1330] & !i[1819]) | ( l_41 [1331] &  i[1819]);
assign l_40[667]    = ( l_41 [1332] & !i[1819]) | ( l_41 [1333] &  i[1819]);
assign l_40[668]    = ( l_41 [1334] & !i[1819]) | ( l_41 [1335] &  i[1819]);
assign l_40[669]    = ( l_41 [1336] & !i[1819]) | ( l_41 [1337] &  i[1819]);
assign l_40[670]    = ( l_41 [1338] & !i[1819]) | ( l_41 [1339] &  i[1819]);
assign l_40[671]    = ( l_41 [1340] & !i[1819]) | ( l_41 [1341] &  i[1819]);
assign l_40[672]    = ( l_41 [1342] & !i[1819]) | ( l_41 [1343] &  i[1819]);
assign l_40[673]    = ( l_41 [1344] & !i[1819]) | ( l_41 [1345] &  i[1819]);
assign l_40[674]    = ( l_41 [1346] & !i[1819]) | ( l_41 [1347] &  i[1819]);
assign l_40[675]    = ( l_41 [1348] & !i[1819]) | ( l_41 [1349] &  i[1819]);
assign l_40[676]    = ( l_41 [1350] & !i[1819]) | ( l_41 [1351] &  i[1819]);
assign l_40[677]    = ( l_41 [1352] & !i[1819]) | ( l_41 [1353] &  i[1819]);
assign l_40[678]    = ( l_41 [1354] & !i[1819]) | ( l_41 [1355] &  i[1819]);
assign l_40[679]    = ( l_41 [1356] & !i[1819]) | ( l_41 [1357] &  i[1819]);
assign l_40[680]    = ( l_41 [1358] & !i[1819]) | ( l_41 [1359] &  i[1819]);
assign l_40[681]    = ( l_41 [1360] & !i[1819]) | ( l_41 [1361] &  i[1819]);
assign l_40[682]    = ( l_41 [1362] & !i[1819]) | ( l_41 [1363] &  i[1819]);
assign l_40[683]    = ( l_41 [1364] & !i[1819]) | ( l_41 [1365] &  i[1819]);
assign l_40[684]    = ( l_41 [1366] & !i[1819]) | ( l_41 [1367] &  i[1819]);
assign l_40[685]    = ( l_41 [1368] & !i[1819]) | ( l_41 [1369] &  i[1819]);
assign l_40[686]    = ( l_41 [1370] & !i[1819]) | ( l_41 [1371] &  i[1819]);
assign l_40[687]    = ( l_41 [1372] & !i[1819]) | ( l_41 [1373] &  i[1819]);
assign l_40[688]    = ( l_41 [1374] & !i[1819]) | ( l_41 [1375] &  i[1819]);
assign l_40[689]    = ( l_41 [1376] & !i[1819]) | ( l_41 [1377] &  i[1819]);
assign l_40[690]    = ( l_41 [1378] & !i[1819]) | ( l_41 [1379] &  i[1819]);
assign l_40[691]    = ( l_41 [1380] & !i[1819]) | ( l_41 [1381] &  i[1819]);
assign l_40[692]    = ( l_41 [1382] & !i[1819]) | ( l_41 [1383] &  i[1819]);
assign l_40[693]    = ( l_41 [1384] & !i[1819]) | ( l_41 [1385] &  i[1819]);
assign l_40[694]    = ( l_41 [1386] & !i[1819]) | ( l_41 [1387] &  i[1819]);
assign l_40[695]    = ( l_41 [1388] & !i[1819]) | ( l_41 [1389] &  i[1819]);
assign l_40[696]    = ( l_41 [1390] & !i[1819]) | ( l_41 [1391] &  i[1819]);
assign l_40[697]    = ( l_41 [1392] & !i[1819]) | ( l_41 [1393] &  i[1819]);
assign l_40[698]    = ( l_41 [1394] & !i[1819]) | ( l_41 [1395] &  i[1819]);
assign l_40[699]    = ( l_41 [1396] & !i[1819]) | ( l_41 [1397] &  i[1819]);
assign l_40[700]    = ( l_41 [1398] & !i[1819]) | ( l_41 [1399] &  i[1819]);
assign l_40[701]    = ( l_41 [1400] & !i[1819]) | ( l_41 [1401] &  i[1819]);
assign l_40[702]    = ( l_41 [1402] & !i[1819]) | ( l_41 [1403] &  i[1819]);
assign l_40[703]    = ( l_41 [1404] & !i[1819]) | ( l_41 [1405] &  i[1819]);
assign l_40[704]    = ( l_41 [1406] & !i[1819]) | ( l_41 [1407] &  i[1819]);
assign l_40[705]    = ( l_41 [1408] & !i[1819]) | ( l_41 [1409] &  i[1819]);
assign l_40[706]    = ( l_41 [1410] & !i[1819]) | ( l_41 [1411] &  i[1819]);
assign l_40[707]    = ( l_41 [1412] & !i[1819]) | ( l_41 [1413] &  i[1819]);
assign l_40[708]    = ( l_41 [1414] & !i[1819]) | ( l_41 [1415] &  i[1819]);
assign l_40[709]    = ( l_41 [1416] & !i[1819]) | ( l_41 [1417] &  i[1819]);
assign l_40[710]    = ( l_41 [1418] & !i[1819]) | ( l_41 [1419] &  i[1819]);
assign l_40[711]    = ( l_41 [1420] & !i[1819]) | ( l_41 [1421] &  i[1819]);
assign l_40[712]    = ( l_41 [1422] & !i[1819]) | ( l_41 [1423] &  i[1819]);
assign l_40[713]    = ( l_41 [1424] & !i[1819]) | ( l_41 [1425] &  i[1819]);
assign l_40[714]    = ( l_41 [1426] & !i[1819]) | ( l_41 [1427] &  i[1819]);
assign l_40[715]    = ( l_41 [1428] & !i[1819]) | ( l_41 [1429] &  i[1819]);
assign l_40[716]    = ( l_41 [1430] & !i[1819]) | ( l_41 [1431] &  i[1819]);
assign l_40[717]    = ( l_41 [1432] & !i[1819]) | ( l_41 [1433] &  i[1819]);
assign l_40[718]    = ( l_41 [1434] & !i[1819]) | ( l_41 [1435] &  i[1819]);
assign l_40[719]    = ( l_41 [1436] & !i[1819]) | ( l_41 [1437] &  i[1819]);
assign l_40[720]    = ( l_41 [1438] & !i[1819]) | ( l_41 [1439] &  i[1819]);
assign l_40[721]    = ( l_41 [1440] & !i[1819]) | ( l_41 [1441] &  i[1819]);
assign l_40[722]    = ( l_41 [1442] & !i[1819]) | ( l_41 [1443] &  i[1819]);
assign l_40[723]    = ( l_41 [1444] & !i[1819]) | ( l_41 [1445] &  i[1819]);
assign l_40[724]    = ( l_41 [1446] & !i[1819]) | ( l_41 [1447] &  i[1819]);
assign l_40[725]    = ( l_41 [1448] & !i[1819]) | ( l_41 [1449] &  i[1819]);
assign l_40[726]    = ( l_41 [1450] & !i[1819]) | ( l_41 [1451] &  i[1819]);
assign l_40[727]    = ( l_41 [1452] & !i[1819]) | ( l_41 [1453] &  i[1819]);
assign l_40[728]    = ( l_41 [1454] & !i[1819]) | ( l_41 [1455] &  i[1819]);
assign l_40[729]    = ( l_41 [1456] & !i[1819]) | ( l_41 [1457] &  i[1819]);
assign l_40[730]    = ( l_41 [1458] & !i[1819]) | ( l_41 [1459] &  i[1819]);
assign l_40[731]    = ( l_41 [1460] & !i[1819]) | ( l_41 [1461] &  i[1819]);
assign l_40[732]    = ( l_41 [1462] & !i[1819]) | ( l_41 [1463] &  i[1819]);
assign l_40[733]    = ( l_41 [1464] & !i[1819]) | ( l_41 [1465] &  i[1819]);
assign l_40[734]    = ( l_41 [1466] & !i[1819]) | ( l_41 [1467] &  i[1819]);
assign l_40[735]    = ( l_41 [1468] & !i[1819]) | ( l_41 [1469] &  i[1819]);
assign l_40[736]    = ( l_41 [1470] & !i[1819]) | ( l_41 [1471] &  i[1819]);
assign l_40[737]    = ( l_41 [1472] & !i[1819]) | ( l_41 [1473] &  i[1819]);
assign l_40[738]    = ( l_41 [1474] & !i[1819]) | ( l_41 [1475] &  i[1819]);
assign l_40[739]    = ( l_41 [1476] & !i[1819]) | ( l_41 [1477] &  i[1819]);
assign l_40[740]    = ( l_41 [1478] & !i[1819]) | ( l_41 [1479] &  i[1819]);
assign l_40[741]    = ( l_41 [1480] & !i[1819]) | ( l_41 [1481] &  i[1819]);
assign l_40[742]    = ( l_41 [1482] & !i[1819]) | ( l_41 [1483] &  i[1819]);
assign l_40[743]    = ( l_41 [1484] & !i[1819]) | ( l_41 [1485] &  i[1819]);
assign l_40[744]    = ( l_41 [1486] & !i[1819]) | ( l_41 [1487] &  i[1819]);
assign l_40[745]    = ( l_41 [1488] & !i[1819]) | ( l_41 [1489] &  i[1819]);
assign l_40[746]    = ( l_41 [1490] & !i[1819]) | ( l_41 [1491] &  i[1819]);
assign l_40[747]    = ( l_41 [1492] & !i[1819]) | ( l_41 [1493] &  i[1819]);
assign l_40[748]    = ( l_41 [1494] & !i[1819]) | ( l_41 [1495] &  i[1819]);
assign l_40[749]    = ( l_41 [1496] & !i[1819]) | ( l_41 [1497] &  i[1819]);
assign l_40[750]    = ( l_41 [1498] & !i[1819]) | ( l_41 [1499] &  i[1819]);
assign l_40[751]    = ( l_41 [1500] & !i[1819]) | ( l_41 [1501] &  i[1819]);
assign l_40[752]    = ( l_41 [1502] & !i[1819]) | ( l_41 [1503] &  i[1819]);
assign l_40[753]    = ( l_41 [1504] & !i[1819]) | ( l_41 [1505] &  i[1819]);
assign l_40[754]    = ( l_41 [1506] & !i[1819]) | ( l_41 [1507] &  i[1819]);
assign l_40[755]    = ( l_41 [1508] & !i[1819]) | ( l_41 [1509] &  i[1819]);
assign l_40[756]    = ( l_41 [1510] & !i[1819]) | ( l_41 [1511] &  i[1819]);
assign l_40[757]    = ( l_41 [1512] & !i[1819]) | ( l_41 [1513] &  i[1819]);
assign l_40[758]    = ( l_41 [1514] & !i[1819]) | ( l_41 [1515] &  i[1819]);
assign l_40[759]    = ( l_41 [1516] & !i[1819]) | ( l_41 [1517] &  i[1819]);
assign l_40[760]    = ( l_41 [1518] & !i[1819]) | ( l_41 [1519] &  i[1819]);
assign l_40[761]    = ( l_41 [1520] & !i[1819]) | ( l_41 [1521] &  i[1819]);
assign l_40[762]    = ( l_41 [1522] & !i[1819]) | ( l_41 [1523] &  i[1819]);
assign l_40[763]    = ( l_41 [1524] & !i[1819]) | ( l_41 [1525] &  i[1819]);
assign l_40[764]    = ( l_41 [1526] & !i[1819]) | ( l_41 [1527] &  i[1819]);
assign l_40[765]    = ( l_41 [1528] & !i[1819]) | ( l_41 [1529] &  i[1819]);
assign l_40[766]    = ( l_41 [1530] & !i[1819]) | ( l_41 [1531] &  i[1819]);
assign l_40[767]    = ( l_41 [1532] & !i[1819]) | ( l_41 [1533] &  i[1819]);
assign l_40[768]    = ( l_41 [1534] & !i[1819]) | ( l_41 [1535] &  i[1819]);
assign l_40[769]    = ( l_41 [1536] & !i[1819]) | ( l_41 [1537] &  i[1819]);
assign l_40[770]    = ( l_41 [1538] & !i[1819]) | ( l_41 [1539] &  i[1819]);
assign l_40[771]    = ( l_41 [1540] & !i[1819]) | ( l_41 [1541] &  i[1819]);
assign l_40[772]    = ( l_41 [1542] & !i[1819]) | ( l_41 [1543] &  i[1819]);
assign l_40[773]    = ( l_41 [1544] & !i[1819]) | ( l_41 [1545] &  i[1819]);
assign l_40[774]    = ( l_41 [1546] & !i[1819]) | ( l_41 [1547] &  i[1819]);
assign l_40[775]    = ( l_41 [1548] & !i[1819]) | ( l_41 [1549] &  i[1819]);
assign l_40[776]    = ( l_41 [1550] & !i[1819]) | ( l_41 [1551] &  i[1819]);
assign l_40[777]    = ( l_41 [1552] & !i[1819]) | ( l_41 [1553] &  i[1819]);
assign l_40[778]    = ( l_41 [1554] & !i[1819]) | ( l_41 [1555] &  i[1819]);
assign l_40[779]    = ( l_41 [1556] & !i[1819]) | ( l_41 [1557] &  i[1819]);
assign l_40[780]    = ( l_41 [1558] & !i[1819]) | ( l_41 [1559] &  i[1819]);
assign l_40[781]    = ( l_41 [1560] & !i[1819]) | ( l_41 [1561] &  i[1819]);
assign l_40[782]    = ( l_41 [1562] & !i[1819]) | ( l_41 [1563] &  i[1819]);
assign l_40[783]    = ( l_41 [1564] & !i[1819]) | ( l_41 [1565] &  i[1819]);
assign l_40[784]    = ( l_41 [1566] & !i[1819]) | ( l_41 [1567] &  i[1819]);
assign l_40[785]    = ( l_41 [1568] & !i[1819]) | ( l_41 [1569] &  i[1819]);
assign l_40[786]    = ( l_41 [1570] & !i[1819]) | ( l_41 [1571] &  i[1819]);
assign l_40[787]    = ( l_41 [1572] & !i[1819]) | ( l_41 [1573] &  i[1819]);
assign l_40[788]    = ( l_41 [1574] & !i[1819]) | ( l_41 [1575] &  i[1819]);
assign l_40[789]    = ( l_41 [1576] & !i[1819]) | ( l_41 [1577] &  i[1819]);
assign l_40[790]    = ( l_41 [1578] & !i[1819]) | ( l_41 [1579] &  i[1819]);
assign l_40[791]    = ( l_41 [1580] & !i[1819]) | ( l_41 [1581] &  i[1819]);
assign l_40[792]    = ( l_41 [1582] & !i[1819]) | ( l_41 [1583] &  i[1819]);
assign l_40[793]    = ( l_41 [1584] & !i[1819]) | ( l_41 [1585] &  i[1819]);
assign l_40[794]    = ( l_41 [1586] & !i[1819]) | ( l_41 [1587] &  i[1819]);
assign l_40[795]    = ( l_41 [1588] & !i[1819]) | ( l_41 [1589] &  i[1819]);
assign l_40[796]    = ( l_41 [1590] & !i[1819]) | ( l_41 [1591] &  i[1819]);
assign l_40[797]    = ( l_41 [1592] & !i[1819]) | ( l_41 [1593] &  i[1819]);
assign l_40[798]    = ( l_41 [1594] & !i[1819]) | ( l_41 [1595] &  i[1819]);
assign l_40[799]    = ( l_41 [1596] & !i[1819]) | ( l_41 [1597] &  i[1819]);
assign l_40[800]    = ( l_41 [1598] & !i[1819]) | ( l_41 [1599] &  i[1819]);
assign l_40[801]    = ( l_41 [1600] & !i[1819]) | ( l_41 [1601] &  i[1819]);
assign l_40[802]    = ( l_41 [1602] & !i[1819]) | ( l_41 [1603] &  i[1819]);
assign l_40[803]    = ( l_41 [1604] & !i[1819]) | ( l_41 [1605] &  i[1819]);
assign l_40[804]    = ( l_41 [1606] & !i[1819]) | ( l_41 [1607] &  i[1819]);
assign l_40[805]    = ( l_41 [1608] & !i[1819]) | ( l_41 [1609] &  i[1819]);
assign l_40[806]    = ( l_41 [1610] & !i[1819]) | ( l_41 [1611] &  i[1819]);
assign l_40[807]    = ( l_41 [1612] & !i[1819]) | ( l_41 [1613] &  i[1819]);
assign l_40[808]    = ( l_41 [1614] & !i[1819]) | ( l_41 [1615] &  i[1819]);
assign l_40[809]    = ( l_41 [1616] & !i[1819]) | ( l_41 [1617] &  i[1819]);
assign l_40[810]    = ( l_41 [1618] & !i[1819]) | ( l_41 [1619] &  i[1819]);
assign l_40[811]    = ( l_41 [1620] & !i[1819]) | ( l_41 [1621] &  i[1819]);
assign l_40[812]    = ( l_41 [1622] & !i[1819]) | ( l_41 [1623] &  i[1819]);
assign l_40[813]    = ( l_41 [1624] & !i[1819]) | ( l_41 [1625] &  i[1819]);
assign l_40[814]    = ( l_41 [1626] & !i[1819]) | ( l_41 [1627] &  i[1819]);
assign l_40[815]    = ( l_41 [1628] & !i[1819]) | ( l_41 [1629] &  i[1819]);
assign l_40[816]    = ( l_41 [1630] & !i[1819]) | ( l_41 [1631] &  i[1819]);
assign l_40[817]    = ( l_41 [1632] & !i[1819]) | ( l_41 [1633] &  i[1819]);
assign l_40[818]    = ( l_41 [1634] & !i[1819]) | ( l_41 [1635] &  i[1819]);
assign l_40[819]    = ( l_41 [1636] & !i[1819]) | ( l_41 [1637] &  i[1819]);
assign l_40[820]    = ( l_41 [1638] & !i[1819]) | ( l_41 [1639] &  i[1819]);
assign l_40[821]    = ( l_41 [1640] & !i[1819]) | ( l_41 [1641] &  i[1819]);
assign l_40[822]    = ( l_41 [1642] & !i[1819]) | ( l_41 [1643] &  i[1819]);
assign l_40[823]    = ( l_41 [1644] & !i[1819]) | ( l_41 [1645] &  i[1819]);
assign l_40[824]    = ( l_41 [1646] & !i[1819]) | ( l_41 [1647] &  i[1819]);
assign l_40[825]    = ( l_41 [1648] & !i[1819]) | ( l_41 [1649] &  i[1819]);
assign l_40[826]    = ( l_41 [1650] & !i[1819]) | ( l_41 [1651] &  i[1819]);
assign l_40[827]    = ( l_41 [1652] & !i[1819]) | ( l_41 [1653] &  i[1819]);
assign l_40[828]    = ( l_41 [1654] & !i[1819]) | ( l_41 [1655] &  i[1819]);
assign l_40[829]    = ( l_41 [1656] & !i[1819]) | ( l_41 [1657] &  i[1819]);
assign l_40[830]    = ( l_41 [1658] & !i[1819]) | ( l_41 [1659] &  i[1819]);
assign l_40[831]    = ( l_41 [1660] & !i[1819]) | ( l_41 [1661] &  i[1819]);
assign l_40[832]    = ( l_41 [1662] & !i[1819]) | ( l_41 [1663] &  i[1819]);
assign l_40[833]    = ( l_41 [1664] & !i[1819]) | ( l_41 [1665] &  i[1819]);
assign l_40[834]    = ( l_41 [1666] & !i[1819]) | ( l_41 [1667] &  i[1819]);
assign l_40[835]    = ( l_41 [1668] & !i[1819]) | ( l_41 [1669] &  i[1819]);
assign l_40[836]    = ( l_41 [1670] & !i[1819]) | ( l_41 [1671] &  i[1819]);
assign l_40[837]    = ( l_41 [1672] & !i[1819]) | ( l_41 [1673] &  i[1819]);
assign l_40[838]    = ( l_41 [1674] & !i[1819]) | ( l_41 [1675] &  i[1819]);
assign l_40[839]    = ( l_41 [1676] & !i[1819]) | ( l_41 [1677] &  i[1819]);
assign l_40[840]    = ( l_41 [1678] & !i[1819]) | ( l_41 [1679] &  i[1819]);
assign l_40[841]    = ( l_41 [1680] & !i[1819]) | ( l_41 [1681] &  i[1819]);
assign l_40[842]    = ( l_41 [1682] & !i[1819]) | ( l_41 [1683] &  i[1819]);
assign l_40[843]    = ( l_41 [1684] & !i[1819]) | ( l_41 [1685] &  i[1819]);
assign l_40[844]    = ( l_41 [1686] & !i[1819]) | ( l_41 [1687] &  i[1819]);
assign l_40[845]    = ( l_41 [1688] & !i[1819]) | ( l_41 [1689] &  i[1819]);
assign l_40[846]    = ( l_41 [1690] & !i[1819]) | ( l_41 [1691] &  i[1819]);
assign l_40[847]    = ( l_41 [1692] & !i[1819]) | ( l_41 [1693] &  i[1819]);
assign l_40[848]    = ( l_41 [1694] & !i[1819]) | ( l_41 [1695] &  i[1819]);
assign l_40[849]    = ( l_41 [1696] & !i[1819]) | ( l_41 [1697] &  i[1819]);
assign l_40[850]    = ( l_41 [1698] & !i[1819]) | ( l_41 [1699] &  i[1819]);
assign l_40[851]    = ( l_41 [1700] & !i[1819]) | ( l_41 [1701] &  i[1819]);
assign l_40[852]    = ( l_41 [1702] & !i[1819]) | ( l_41 [1703] &  i[1819]);
assign l_40[853]    = ( l_41 [1704] & !i[1819]) | ( l_41 [1705] &  i[1819]);
assign l_40[854]    = ( l_41 [1706] & !i[1819]) | ( l_41 [1707] &  i[1819]);
assign l_40[855]    = ( l_41 [1708] & !i[1819]) | ( l_41 [1709] &  i[1819]);
assign l_40[856]    = ( l_41 [1710] & !i[1819]) | ( l_41 [1711] &  i[1819]);
assign l_40[857]    = ( l_41 [1712] & !i[1819]) | ( l_41 [1713] &  i[1819]);
assign l_40[858]    = ( l_41 [1714] & !i[1819]) | ( l_41 [1715] &  i[1819]);
assign l_40[859]    = ( l_41 [1716] & !i[1819]) | ( l_41 [1717] &  i[1819]);
assign l_40[860]    = ( l_41 [1718] & !i[1819]) | ( l_41 [1719] &  i[1819]);
assign l_40[861]    = ( l_41 [1720] & !i[1819]) | ( l_41 [1721] &  i[1819]);
assign l_40[862]    = ( l_41 [1722] & !i[1819]) | ( l_41 [1723] &  i[1819]);
assign l_40[863]    = ( l_41 [1724] & !i[1819]) | ( l_41 [1725] &  i[1819]);
assign l_40[864]    = ( l_41 [1726] & !i[1819]) | ( l_41 [1727] &  i[1819]);
assign l_40[865]    = ( l_41 [1728] & !i[1819]) | ( l_41 [1729] &  i[1819]);
assign l_40[866]    = ( l_41 [1730] & !i[1819]) | ( l_41 [1731] &  i[1819]);
assign l_40[867]    = ( l_41 [1732] & !i[1819]) | ( l_41 [1733] &  i[1819]);
assign l_40[868]    = ( l_41 [1734] & !i[1819]) | ( l_41 [1735] &  i[1819]);
assign l_40[869]    = ( l_41 [1736] & !i[1819]) | ( l_41 [1737] &  i[1819]);
assign l_40[870]    = ( l_41 [1738] & !i[1819]) | ( l_41 [1739] &  i[1819]);
assign l_40[871]    = ( l_41 [1740] & !i[1819]) | ( l_41 [1741] &  i[1819]);
assign l_40[872]    = ( l_41 [1742] & !i[1819]) | ( l_41 [1743] &  i[1819]);
assign l_40[873]    = ( l_41 [1744] & !i[1819]) | ( l_41 [1745] &  i[1819]);
assign l_40[874]    = ( l_41 [1746] & !i[1819]) | ( l_41 [1747] &  i[1819]);
assign l_40[875]    = ( l_41 [1748] & !i[1819]) | ( l_41 [1749] &  i[1819]);
assign l_40[876]    = ( l_41 [1750] & !i[1819]) | ( l_41 [1751] &  i[1819]);
assign l_40[877]    = ( l_41 [1752] & !i[1819]) | ( l_41 [1753] &  i[1819]);
assign l_40[878]    = ( l_41 [1754] & !i[1819]) | ( l_41 [1755] &  i[1819]);
assign l_40[879]    = ( l_41 [1756] & !i[1819]) | ( l_41 [1757] &  i[1819]);
assign l_40[880]    = ( l_41 [1758] & !i[1819]) | ( l_41 [1759] &  i[1819]);
assign l_40[881]    = ( l_41 [1760] & !i[1819]) | ( l_41 [1761] &  i[1819]);
assign l_40[882]    = ( l_41 [1762] & !i[1819]) | ( l_41 [1763] &  i[1819]);
assign l_40[883]    = ( l_41 [1764] & !i[1819]) | ( l_41 [1765] &  i[1819]);
assign l_40[884]    = ( l_41 [1766] & !i[1819]) | ( l_41 [1767] &  i[1819]);
assign l_40[885]    = ( l_41 [1768] & !i[1819]) | ( l_41 [1769] &  i[1819]);
assign l_40[886]    = ( l_41 [1770] & !i[1819]) | ( l_41 [1771] &  i[1819]);
assign l_40[887]    = ( l_41 [1772] & !i[1819]) | ( l_41 [1773] &  i[1819]);
assign l_40[888]    = ( l_41 [1774] & !i[1819]) | ( l_41 [1775] &  i[1819]);
assign l_40[889]    = ( l_41 [1776] & !i[1819]) | ( l_41 [1777] &  i[1819]);
assign l_40[890]    = ( l_41 [1778] & !i[1819]) | ( l_41 [1779] &  i[1819]);
assign l_40[891]    = ( l_41 [1780] & !i[1819]) | ( l_41 [1781] &  i[1819]);
assign l_40[892]    = ( l_41 [1782] & !i[1819]) | ( l_41 [1783] &  i[1819]);
assign l_40[893]    = ( l_41 [1784] & !i[1819]) | ( l_41 [1785] &  i[1819]);
assign l_40[894]    = ( l_41 [1786] & !i[1819]) | ( l_41 [1787] &  i[1819]);
assign l_40[895]    = ( l_41 [1788] & !i[1819]) | ( l_41 [1789] &  i[1819]);
assign l_40[896]    = ( l_41 [1790] & !i[1819]) | ( l_41 [1791] &  i[1819]);
assign l_40[897]    = ( l_41 [1792] & !i[1819]) | ( l_41 [1793] &  i[1819]);
assign l_40[898]    = ( l_41 [1794] & !i[1819]) | ( l_41 [1795] &  i[1819]);
assign l_40[899]    = ( l_41 [1796] & !i[1819]) | ( l_41 [1797] &  i[1819]);
assign l_40[900]    = ( l_41 [1798] & !i[1819]) | ( l_41 [1799] &  i[1819]);
assign l_40[901]    = ( l_41 [1800] & !i[1819]) | ( l_41 [1801] &  i[1819]);
assign l_40[902]    = ( l_41 [1802] & !i[1819]) | ( l_41 [1803] &  i[1819]);
assign l_40[903]    = ( l_41 [1804] & !i[1819]) | ( l_41 [1805] &  i[1819]);
assign l_40[904]    = ( l_41 [1806] & !i[1819]) | ( l_41 [1807] &  i[1819]);
assign l_40[905]    = ( l_41 [1808] & !i[1819]) | ( l_41 [1809] &  i[1819]);
assign l_40[906]    = ( l_41 [1810] & !i[1819]) | ( l_41 [1811] &  i[1819]);
assign l_40[907]    = ( l_41 [1812] & !i[1819]) | ( l_41 [1813] &  i[1819]);
assign l_40[908]    = ( l_41 [1814] & !i[1819]) | ( l_41 [1815] &  i[1819]);
assign l_40[909]    = ( l_41 [1816] & !i[1819]) | ( l_41 [1817] &  i[1819]);
assign l_40[910]    = ( l_41 [1818] & !i[1819]) | ( l_41 [1819] &  i[1819]);
assign l_40[911]    = ( l_41 [1820] & !i[1819]) | ( l_41 [1821] &  i[1819]);
assign l_40[912]    = ( l_41 [1822] & !i[1819]) | ( l_41 [1823] &  i[1819]);
assign l_40[913]    = ( l_41 [1824] & !i[1819]) | ( l_41 [1825] &  i[1819]);
assign l_40[914]    = ( l_41 [1826] & !i[1819]) | ( l_41 [1827] &  i[1819]);
assign l_40[915]    = ( l_41 [1828] & !i[1819]) | ( l_41 [1829] &  i[1819]);
assign l_40[916]    = ( l_41 [1830] & !i[1819]) | ( l_41 [1831] &  i[1819]);
assign l_40[917]    = ( l_41 [1832] & !i[1819]) | ( l_41 [1833] &  i[1819]);
assign l_40[918]    = ( l_41 [1834] & !i[1819]) | ( l_41 [1835] &  i[1819]);
assign l_40[919]    = ( l_41 [1836] & !i[1819]) | ( l_41 [1837] &  i[1819]);
assign l_40[920]    = ( l_41 [1838] & !i[1819]) | ( l_41 [1839] &  i[1819]);
assign l_40[921]    = ( l_41 [1840] & !i[1819]) | ( l_41 [1841] &  i[1819]);
assign l_40[922]    = ( l_41 [1842] & !i[1819]) | ( l_41 [1843] &  i[1819]);
assign l_40[923]    = ( l_41 [1844] & !i[1819]) | ( l_41 [1845] &  i[1819]);
assign l_40[924]    = ( l_41 [1846] & !i[1819]) | ( l_41 [1847] &  i[1819]);
assign l_40[925]    = ( l_41 [1848] & !i[1819]) | ( l_41 [1849] &  i[1819]);
assign l_40[926]    = ( l_41 [1850] & !i[1819]) | ( l_41 [1851] &  i[1819]);
assign l_40[927]    = ( l_41 [1852] & !i[1819]) | ( l_41 [1853] &  i[1819]);
assign l_40[928]    = ( l_41 [1854] & !i[1819]) | ( l_41 [1855] &  i[1819]);
assign l_40[929]    = ( l_41 [1856] & !i[1819]) | ( l_41 [1857] &  i[1819]);
assign l_40[930]    = ( l_41 [1858] & !i[1819]) | ( l_41 [1859] &  i[1819]);
assign l_40[931]    = ( l_41 [1860] & !i[1819]) | ( l_41 [1861] &  i[1819]);
assign l_40[932]    = ( l_41 [1862] & !i[1819]) | ( l_41 [1863] &  i[1819]);
assign l_40[933]    = ( l_41 [1864] & !i[1819]) | ( l_41 [1865] &  i[1819]);
assign l_40[934]    = ( l_41 [1866] & !i[1819]) | ( l_41 [1867] &  i[1819]);
assign l_40[935]    = ( l_41 [1868] & !i[1819]) | ( l_41 [1869] &  i[1819]);
assign l_40[936]    = ( l_41 [1870] & !i[1819]) | ( l_41 [1871] &  i[1819]);
assign l_40[937]    = ( l_41 [1872] & !i[1819]) | ( l_41 [1873] &  i[1819]);
assign l_40[938]    = ( l_41 [1874] & !i[1819]) | ( l_41 [1875] &  i[1819]);
assign l_40[939]    = ( l_41 [1876] & !i[1819]) | ( l_41 [1877] &  i[1819]);
assign l_40[940]    = ( l_41 [1878] & !i[1819]) | ( l_41 [1879] &  i[1819]);
assign l_40[941]    = ( l_41 [1880] & !i[1819]) | ( l_41 [1881] &  i[1819]);
assign l_40[942]    = ( l_41 [1882] & !i[1819]) | ( l_41 [1883] &  i[1819]);
assign l_40[943]    = ( l_41 [1884] & !i[1819]) | ( l_41 [1885] &  i[1819]);
assign l_40[944]    = ( l_41 [1886] & !i[1819]) | ( l_41 [1887] &  i[1819]);
assign l_40[945]    = ( l_41 [1888] & !i[1819]) | ( l_41 [1889] &  i[1819]);
assign l_40[946]    = ( l_41 [1890] & !i[1819]) | ( l_41 [1891] &  i[1819]);
assign l_40[947]    = ( l_41 [1892] & !i[1819]) | ( l_41 [1893] &  i[1819]);
assign l_40[948]    = ( l_41 [1894] & !i[1819]) | ( l_41 [1895] &  i[1819]);
assign l_40[949]    = ( l_41 [1896] & !i[1819]) | ( l_41 [1897] &  i[1819]);
assign l_40[950]    = ( l_41 [1898] & !i[1819]) | ( l_41 [1899] &  i[1819]);
assign l_40[951]    = ( l_41 [1900] & !i[1819]) | ( l_41 [1901] &  i[1819]);
assign l_40[952]    = ( l_41 [1902] & !i[1819]) | ( l_41 [1903] &  i[1819]);
assign l_40[953]    = ( l_41 [1904] & !i[1819]) | ( l_41 [1905] &  i[1819]);
assign l_40[954]    = ( l_41 [1906] & !i[1819]) | ( l_41 [1907] &  i[1819]);
assign l_40[955]    = ( l_41 [1908] & !i[1819]) | ( l_41 [1909] &  i[1819]);
assign l_40[956]    = ( l_41 [1910] & !i[1819]) | ( l_41 [1911] &  i[1819]);
assign l_40[957]    = ( l_41 [1912] & !i[1819]) | ( l_41 [1913] &  i[1819]);
assign l_40[958]    = ( l_41 [1914] & !i[1819]) | ( l_41 [1915] &  i[1819]);
assign l_40[959]    = ( l_41 [1916] & !i[1819]) | ( l_41 [1917] &  i[1819]);
assign l_40[960]    = ( l_41 [1918] & !i[1819]) | ( l_41 [1919] &  i[1819]);
assign l_40[961]    = ( l_41 [1920] & !i[1819]) | ( l_41 [1921] &  i[1819]);
assign l_40[962]    = ( l_41 [1922] & !i[1819]) | ( l_41 [1923] &  i[1819]);
assign l_40[963]    = ( l_41 [1924] & !i[1819]) | ( l_41 [1925] &  i[1819]);
assign l_40[964]    = ( l_41 [1926] & !i[1819]) | ( l_41 [1927] &  i[1819]);
assign l_40[965]    = ( l_41 [1928] & !i[1819]) | ( l_41 [1929] &  i[1819]);
assign l_40[966]    = ( l_41 [1930] & !i[1819]) | ( l_41 [1931] &  i[1819]);
assign l_40[967]    = ( l_41 [1932] & !i[1819]) | ( l_41 [1933] &  i[1819]);
assign l_40[968]    = ( l_41 [1934] & !i[1819]) | ( l_41 [1935] &  i[1819]);
assign l_40[969]    = ( l_41 [1936] & !i[1819]) | ( l_41 [1937] &  i[1819]);
assign l_40[970]    = ( l_41 [1938] & !i[1819]) | ( l_41 [1939] &  i[1819]);
assign l_40[971]    = ( l_41 [1940] & !i[1819]) | ( l_41 [1941] &  i[1819]);
assign l_40[972]    = ( l_41 [1942] & !i[1819]) | ( l_41 [1943] &  i[1819]);
assign l_40[973]    = ( l_41 [1944] & !i[1819]) | ( l_41 [1945] &  i[1819]);
assign l_40[974]    = ( l_41 [1946] & !i[1819]) | ( l_41 [1947] &  i[1819]);
assign l_40[975]    = ( l_41 [1948] & !i[1819]) | ( l_41 [1949] &  i[1819]);
assign l_40[976]    = ( l_41 [1950] & !i[1819]) | ( l_41 [1951] &  i[1819]);
assign l_40[977]    = ( l_41 [1952] & !i[1819]) | ( l_41 [1953] &  i[1819]);
assign l_40[978]    = ( l_41 [1954] & !i[1819]) | ( l_41 [1955] &  i[1819]);
assign l_40[979]    = ( l_41 [1956] & !i[1819]) | ( l_41 [1957] &  i[1819]);
assign l_40[980]    = ( l_41 [1958] & !i[1819]) | ( l_41 [1959] &  i[1819]);
assign l_40[981]    = ( l_41 [1960] & !i[1819]) | ( l_41 [1961] &  i[1819]);
assign l_40[982]    = ( l_41 [1962] & !i[1819]) | ( l_41 [1963] &  i[1819]);
assign l_40[983]    = ( l_41 [1964] & !i[1819]) | ( l_41 [1965] &  i[1819]);
assign l_40[984]    = ( l_41 [1966] & !i[1819]) | ( l_41 [1967] &  i[1819]);
assign l_40[985]    = ( l_41 [1968] & !i[1819]) | ( l_41 [1969] &  i[1819]);
assign l_40[986]    = ( l_41 [1970] & !i[1819]) | ( l_41 [1971] &  i[1819]);
assign l_40[987]    = ( l_41 [1972] & !i[1819]) | ( l_41 [1973] &  i[1819]);
assign l_40[988]    = ( l_41 [1974] & !i[1819]) | ( l_41 [1975] &  i[1819]);
assign l_40[989]    = ( l_41 [1976] & !i[1819]) | ( l_41 [1977] &  i[1819]);
assign l_40[990]    = ( l_41 [1978] & !i[1819]) | ( l_41 [1979] &  i[1819]);
assign l_40[991]    = ( l_41 [1980] & !i[1819]) | ( l_41 [1981] &  i[1819]);
assign l_40[992]    = ( l_41 [1982] & !i[1819]) | ( l_41 [1983] &  i[1819]);
assign l_40[993]    = ( l_41 [1984] & !i[1819]) | ( l_41 [1985] &  i[1819]);
assign l_40[994]    = ( l_41 [1986] & !i[1819]) | ( l_41 [1987] &  i[1819]);
assign l_40[995]    = ( l_41 [1988] & !i[1819]) | ( l_41 [1989] &  i[1819]);
assign l_40[996]    = ( l_41 [1990] & !i[1819]) | ( l_41 [1991] &  i[1819]);
assign l_40[997]    = ( l_41 [1992] & !i[1819]) | ( l_41 [1993] &  i[1819]);
assign l_40[998]    = ( l_41 [1994] & !i[1819]) | ( l_41 [1995] &  i[1819]);
assign l_40[999]    = ( l_41 [1996] & !i[1819]) | ( l_41 [1997] &  i[1819]);
assign l_40[1000]    = ( l_41 [1998] & !i[1819]) | ( l_41 [1999] &  i[1819]);
assign l_40[1001]    = ( l_41 [2000] & !i[1819]) | ( l_41 [2001] &  i[1819]);
assign l_40[1002]    = ( l_41 [2002] & !i[1819]) | ( l_41 [2003] &  i[1819]);
assign l_40[1003]    = ( l_41 [2004] & !i[1819]) | ( l_41 [2005] &  i[1819]);
assign l_40[1004]    = ( l_41 [2006] & !i[1819]) | ( l_41 [2007] &  i[1819]);
assign l_40[1005]    = ( l_41 [2008] & !i[1819]) | ( l_41 [2009] &  i[1819]);
assign l_40[1006]    = ( l_41 [2010] & !i[1819]) | ( l_41 [2011] &  i[1819]);
assign l_40[1007]    = ( l_41 [2012] & !i[1819]) | ( l_41 [2013] &  i[1819]);
assign l_40[1008]    = ( l_41 [2014] & !i[1819]) | ( l_41 [2015] &  i[1819]);
assign l_40[1009]    = ( l_41 [2016] & !i[1819]) | ( l_41 [2017] &  i[1819]);
assign l_40[1010]    = ( l_41 [2018] & !i[1819]) | ( l_41 [2019] &  i[1819]);
assign l_40[1011]    = ( l_41 [2020] & !i[1819]) | ( l_41 [2021] &  i[1819]);
assign l_40[1012]    = ( l_41 [2022] & !i[1819]) | ( l_41 [2023] &  i[1819]);
assign l_40[1013]    = ( l_41 [2024] & !i[1819]) | ( l_41 [2025] &  i[1819]);
assign l_40[1014]    = ( l_41 [2026] & !i[1819]) | ( l_41 [2027] &  i[1819]);
assign l_40[1015]    = ( l_41 [2028] & !i[1819]) | ( l_41 [2029] &  i[1819]);
assign l_40[1016]    = ( l_41 [2030] & !i[1819]) | ( l_41 [2031] &  i[1819]);
assign l_40[1017]    = ( l_41 [2032] & !i[1819]) | ( l_41 [2033] &  i[1819]);
assign l_40[1018]    = ( l_41 [2034] & !i[1819]) | ( l_41 [2035] &  i[1819]);
assign l_40[1019]    = ( l_41 [2036] & !i[1819]) | ( l_41 [2037] &  i[1819]);
assign l_40[1020]    = ( l_41 [2038] & !i[1819]) | ( l_41 [2039] &  i[1819]);
assign l_40[1021]    = ( l_41 [2040] & !i[1819]) | ( l_41 [2041] &  i[1819]);
assign l_40[1022]    = ( l_41 [2042] & !i[1819]) | ( l_41 [2043] &  i[1819]);
assign l_40[1023]    = ( l_41 [2044] & !i[1819]) | ( l_41 [2045] &  i[1819]);
assign l_40[1024]    = ( l_41 [2046] & !i[1819]) | ( l_41 [2047] &  i[1819]);
assign l_40[1025]    = ( l_41 [2048] & !i[1819]) | ( l_41 [2049] &  i[1819]);
assign l_40[1026]    = ( l_41 [2050] & !i[1819]) | ( l_41 [2051] &  i[1819]);
assign l_40[1027]    = ( l_41 [2052] & !i[1819]) | ( l_41 [2053] &  i[1819]);
assign l_40[1028]    = ( l_41 [2054] & !i[1819]) | ( l_41 [2055] &  i[1819]);
assign l_40[1029]    = ( l_41 [2056] & !i[1819]) | ( l_41 [2057] &  i[1819]);
assign l_40[1030]    = ( l_41 [2058] & !i[1819]) | ( l_41 [2059] &  i[1819]);
assign l_40[1031]    = ( l_41 [2060] & !i[1819]) | ( l_41 [2061] &  i[1819]);
assign l_40[1032]    = ( l_41 [2062] & !i[1819]) | ( l_41 [2063] &  i[1819]);
assign l_40[1033]    = ( l_41 [2064] & !i[1819]) | ( l_41 [2065] &  i[1819]);
assign l_40[1034]    = ( l_41 [2066] & !i[1819]) | ( l_41 [2067] &  i[1819]);
assign l_40[1035]    = ( l_41 [2068] & !i[1819]) | ( l_41 [2069] &  i[1819]);
assign l_40[1036]    = ( l_41 [2070] & !i[1819]) | ( l_41 [2071] &  i[1819]);
assign l_40[1037]    = ( l_41 [2072] & !i[1819]) | ( l_41 [2073] &  i[1819]);
assign l_40[1038]    = ( l_41 [2074] & !i[1819]) | ( l_41 [2075] &  i[1819]);
assign l_40[1039]    = ( l_41 [2076] & !i[1819]) | ( l_41 [2077] &  i[1819]);
assign l_40[1040]    = ( l_41 [2078] & !i[1819]) | ( l_41 [2079] &  i[1819]);
assign l_40[1041]    = ( l_41 [2080] & !i[1819]) | ( l_41 [2081] &  i[1819]);
assign l_40[1042]    = ( l_41 [2082] & !i[1819]) | ( l_41 [2083] &  i[1819]);
assign l_40[1043]    = ( l_41 [2084] & !i[1819]) | ( l_41 [2085] &  i[1819]);
assign l_40[1044]    = ( l_41 [2086] & !i[1819]) | ( l_41 [2087] &  i[1819]);
assign l_40[1045]    = ( l_41 [2088] & !i[1819]) | ( l_41 [2089] &  i[1819]);
assign l_40[1046]    = ( l_41 [2090] & !i[1819]) | ( l_41 [2091] &  i[1819]);
assign l_40[1047]    = ( l_41 [2092] & !i[1819]) | ( l_41 [2093] &  i[1819]);
assign l_40[1048]    = ( l_41 [2094] & !i[1819]) | ( l_41 [2095] &  i[1819]);
assign l_40[1049]    = ( l_41 [2096] & !i[1819]) | ( l_41 [2097] &  i[1819]);
assign l_40[1050]    = ( l_41 [2098] & !i[1819]) | ( l_41 [2099] &  i[1819]);
assign l_40[1051]    = ( l_41 [2100] & !i[1819]) | ( l_41 [2101] &  i[1819]);
assign l_40[1052]    = ( l_41 [2102] & !i[1819]) | ( l_41 [2103] &  i[1819]);
assign l_40[1053]    = ( l_41 [2104] & !i[1819]) | ( l_41 [2105] &  i[1819]);
assign l_40[1054]    = ( l_41 [2106] & !i[1819]) | ( l_41 [2107] &  i[1819]);
assign l_40[1055]    = ( l_41 [2108] & !i[1819]) | ( l_41 [2109] &  i[1819]);
assign l_40[1056]    = ( l_41 [2110] & !i[1819]) | ( l_41 [2111] &  i[1819]);
assign l_40[1057]    = ( l_41 [2112] & !i[1819]) | ( l_41 [2113] &  i[1819]);
assign l_40[1058]    = ( l_41 [2114] & !i[1819]) | ( l_41 [2115] &  i[1819]);
assign l_40[1059]    = ( l_41 [2116] & !i[1819]) | ( l_41 [2117] &  i[1819]);
assign l_40[1060]    = ( l_41 [2118] & !i[1819]) | ( l_41 [2119] &  i[1819]);
assign l_40[1061]    = ( l_41 [2120] & !i[1819]) | ( l_41 [2121] &  i[1819]);
assign l_40[1062]    = ( l_41 [2122] & !i[1819]) | ( l_41 [2123] &  i[1819]);
assign l_40[1063]    = ( l_41 [2124] & !i[1819]) | ( l_41 [2125] &  i[1819]);
assign l_40[1064]    = ( l_41 [2126] & !i[1819]) | ( l_41 [2127] &  i[1819]);
assign l_40[1065]    = ( l_41 [2128] & !i[1819]) | ( l_41 [2129] &  i[1819]);
assign l_40[1066]    = ( l_41 [2130] & !i[1819]) | ( l_41 [2131] &  i[1819]);
assign l_40[1067]    = ( l_41 [2132] & !i[1819]) | ( l_41 [2133] &  i[1819]);
assign l_40[1068]    = ( l_41 [2134] & !i[1819]) | ( l_41 [2135] &  i[1819]);
assign l_40[1069]    = ( l_41 [2136] & !i[1819]) | ( l_41 [2137] &  i[1819]);
assign l_40[1070]    = ( l_41 [2138] & !i[1819]) | ( l_41 [2139] &  i[1819]);
assign l_40[1071]    = ( l_41 [2140] & !i[1819]) | ( l_41 [2141] &  i[1819]);
assign l_40[1072]    = ( l_41 [2142] & !i[1819]) | ( l_41 [2143] &  i[1819]);
assign l_40[1073]    = ( l_41 [2144] & !i[1819]) | ( l_41 [2145] &  i[1819]);
assign l_40[1074]    = ( l_41 [2146] & !i[1819]) | ( l_41 [2147] &  i[1819]);
assign l_40[1075]    = ( l_41 [2148] & !i[1819]) | ( l_41 [2149] &  i[1819]);
assign l_40[1076]    = ( l_41 [2150] & !i[1819]) | ( l_41 [2151] &  i[1819]);
assign l_40[1077]    = ( l_41 [2152] & !i[1819]) | ( l_41 [2153] &  i[1819]);
assign l_40[1078]    = ( l_41 [2154] & !i[1819]) | ( l_41 [2155] &  i[1819]);
assign l_40[1079]    = ( l_41 [2156] & !i[1819]) | ( l_41 [2157] &  i[1819]);
assign l_40[1080]    = ( l_41 [2158] & !i[1819]) | ( l_41 [2159] &  i[1819]);
assign l_40[1081]    = ( l_41 [2160] & !i[1819]) | ( l_41 [2161] &  i[1819]);
assign l_40[1082]    = ( l_41 [2162] & !i[1819]) | ( l_41 [2163] &  i[1819]);
assign l_40[1083]    = ( l_41 [2164] & !i[1819]) | ( l_41 [2165] &  i[1819]);
assign l_40[1084]    = ( l_41 [2166] & !i[1819]) | ( l_41 [2167] &  i[1819]);
assign l_40[1085]    = ( l_41 [2168] & !i[1819]) | ( l_41 [2169] &  i[1819]);
assign l_40[1086]    = ( l_41 [2170] & !i[1819]) | ( l_41 [2171] &  i[1819]);
assign l_40[1087]    = ( l_41 [2172] & !i[1819]) | ( l_41 [2173] &  i[1819]);
assign l_40[1088]    = ( l_41 [2174] & !i[1819]) | ( l_41 [2175] &  i[1819]);
assign l_40[1089]    = ( l_41 [2176] & !i[1819]) | ( l_41 [2177] &  i[1819]);
assign l_40[1090]    = ( l_41 [2178] & !i[1819]) | ( l_41 [2179] &  i[1819]);
assign l_40[1091]    = ( l_41 [2180] & !i[1819]) | ( l_41 [2181] &  i[1819]);
assign l_40[1092]    = ( l_41 [2182] & !i[1819]) | ( l_41 [2183] &  i[1819]);
assign l_40[1093]    = ( l_41 [2184] & !i[1819]) | ( l_41 [2185] &  i[1819]);
assign l_40[1094]    = ( l_41 [2186] & !i[1819]) | ( l_41 [2187] &  i[1819]);
assign l_40[1095]    = ( l_41 [2188] & !i[1819]) | ( l_41 [2189] &  i[1819]);
assign l_40[1096]    = ( l_41 [2190] & !i[1819]) | ( l_41 [2191] &  i[1819]);
assign l_40[1097]    = ( l_41 [2192] & !i[1819]) | ( l_41 [2193] &  i[1819]);
assign l_40[1098]    = ( l_41 [2194] & !i[1819]) | ( l_41 [2195] &  i[1819]);
assign l_40[1099]    = ( l_41 [2196] & !i[1819]) | ( l_41 [2197] &  i[1819]);
assign l_40[1100]    = ( l_41 [2198] & !i[1819]) | ( l_41 [2199] &  i[1819]);
assign l_40[1101]    = ( l_41 [2200] & !i[1819]) | ( l_41 [2201] &  i[1819]);
assign l_40[1102]    = ( l_41 [2202] & !i[1819]) | ( l_41 [2203] &  i[1819]);
assign l_40[1103]    = ( l_41 [2204] & !i[1819]) | ( l_41 [2205] &  i[1819]);
assign l_40[1104]    = ( l_41 [2206] & !i[1819]) | ( l_41 [2207] &  i[1819]);
assign l_40[1105]    = ( l_41 [2208] & !i[1819]) | ( l_41 [2209] &  i[1819]);
assign l_40[1106]    = ( l_41 [2210] & !i[1819]) | ( l_41 [2211] &  i[1819]);
assign l_40[1107]    = ( l_41 [2212] & !i[1819]) | ( l_41 [2213] &  i[1819]);
assign l_40[1108]    = ( l_41 [2214] & !i[1819]) | ( l_41 [2215] &  i[1819]);
assign l_40[1109]    = ( l_41 [2216] & !i[1819]) | ( l_41 [2217] &  i[1819]);
assign l_40[1110]    = ( l_41 [2218] & !i[1819]) | ( l_41 [2219] &  i[1819]);
assign l_40[1111]    = ( l_41 [2220] & !i[1819]) | ( l_41 [2221] &  i[1819]);
assign l_40[1112]    = ( l_41 [2222] & !i[1819]) | ( l_41 [2223] &  i[1819]);
assign l_40[1113]    = ( l_41 [2224] & !i[1819]) | ( l_41 [2225] &  i[1819]);
assign l_40[1114]    = ( l_41 [2226] & !i[1819]) | ( l_41 [2227] &  i[1819]);
assign l_40[1115]    = ( l_41 [2228] & !i[1819]) | ( l_41 [2229] &  i[1819]);
assign l_40[1116]    = ( l_41 [2230] & !i[1819]) | ( l_41 [2231] &  i[1819]);
assign l_40[1117]    = ( l_41 [2232] & !i[1819]) | ( l_41 [2233] &  i[1819]);
assign l_40[1118]    = ( l_41 [2234] & !i[1819]) | ( l_41 [2235] &  i[1819]);
assign l_40[1119]    = ( l_41 [2236] & !i[1819]) | ( l_41 [2237] &  i[1819]);
assign l_40[1120]    = ( l_41 [2238] & !i[1819]) | ( l_41 [2239] &  i[1819]);
assign l_40[1121]    = ( l_41 [2240] & !i[1819]) | ( l_41 [2241] &  i[1819]);
assign l_40[1122]    = ( l_41 [2242] & !i[1819]) | ( l_41 [2243] &  i[1819]);
assign l_40[1123]    = ( l_41 [2244] & !i[1819]) | ( l_41 [2245] &  i[1819]);
assign l_40[1124]    = ( l_41 [2246] & !i[1819]) | ( l_41 [2247] &  i[1819]);
assign l_40[1125]    = ( l_41 [2248] & !i[1819]) | ( l_41 [2249] &  i[1819]);
assign l_40[1126]    = ( l_41 [2250] & !i[1819]) | ( l_41 [2251] &  i[1819]);
assign l_40[1127]    = ( l_41 [2252] & !i[1819]) | ( l_41 [2253] &  i[1819]);
assign l_40[1128]    = ( l_41 [2254] & !i[1819]) | ( l_41 [2255] &  i[1819]);
assign l_40[1129]    = ( l_41 [2256] & !i[1819]) | ( l_41 [2257] &  i[1819]);
assign l_40[1130]    = ( l_41 [2258] & !i[1819]) | ( l_41 [2259] &  i[1819]);
assign l_40[1131]    = ( l_41 [2260] & !i[1819]) | ( l_41 [2261] &  i[1819]);
assign l_40[1132]    = ( l_41 [2262] & !i[1819]) | ( l_41 [2263] &  i[1819]);
assign l_40[1133]    = ( l_41 [2264] & !i[1819]) | ( l_41 [2265] &  i[1819]);
assign l_40[1134]    = ( l_41 [2266] & !i[1819]) | ( l_41 [2267] &  i[1819]);
assign l_40[1135]    = ( l_41 [2268] & !i[1819]) | ( l_41 [2269] &  i[1819]);
assign l_40[1136]    = ( l_41 [2270] & !i[1819]) | ( l_41 [2271] &  i[1819]);
assign l_40[1137]    = ( l_41 [2272] & !i[1819]) | ( l_41 [2273] &  i[1819]);
assign l_40[1138]    = ( l_41 [2274] & !i[1819]) | ( l_41 [2275] &  i[1819]);
assign l_40[1139]    = ( l_41 [2276] & !i[1819]) | ( l_41 [2277] &  i[1819]);
assign l_40[1140]    = ( l_41 [2278] & !i[1819]) | ( l_41 [2279] &  i[1819]);
assign l_40[1141]    = ( l_41 [2280] & !i[1819]) | ( l_41 [2281] &  i[1819]);
assign l_40[1142]    = ( l_41 [2282] & !i[1819]) | ( l_41 [2283] &  i[1819]);
assign l_40[1143]    = ( l_41 [2284] & !i[1819]) | ( l_41 [2285] &  i[1819]);
assign l_40[1144]    = ( l_41 [2286] & !i[1819]) | ( l_41 [2287] &  i[1819]);
assign l_40[1145]    = ( l_41 [2288] & !i[1819]) | ( l_41 [2289] &  i[1819]);
assign l_40[1146]    = ( l_41 [2290] & !i[1819]) | ( l_41 [2291] &  i[1819]);
assign l_40[1147]    = ( l_41 [2292] & !i[1819]) | ( l_41 [2293] &  i[1819]);
assign l_40[1148]    = ( l_41 [2294] & !i[1819]) | ( l_41 [2295] &  i[1819]);
assign l_40[1149]    = ( l_41 [2296] & !i[1819]) | ( l_41 [2297] &  i[1819]);
assign l_40[1150]    = ( l_41 [2298] & !i[1819]) | ( l_41 [2299] &  i[1819]);
assign l_40[1151]    = ( l_41 [2300] & !i[1819]) | ( l_41 [2301] &  i[1819]);
assign l_40[1152]    = ( l_41 [2302] & !i[1819]) | ( l_41 [2303] &  i[1819]);
assign l_40[1153]    = ( l_41 [2304] & !i[1819]) | ( l_41 [2305] &  i[1819]);
assign l_40[1154]    = ( l_41 [2306] & !i[1819]) | ( l_41 [2307] &  i[1819]);
assign l_40[1155]    = ( l_41 [2308] & !i[1819]) | ( l_41 [2309] &  i[1819]);
assign l_40[1156]    = ( l_41 [2310] & !i[1819]) | ( l_41 [2311] &  i[1819]);
assign l_40[1157]    = ( l_41 [2312] & !i[1819]) | ( l_41 [2313] &  i[1819]);
assign l_40[1158]    = ( l_41 [2314] & !i[1819]) | ( l_41 [2315] &  i[1819]);
assign l_40[1159]    = ( l_41 [2316] & !i[1819]) | ( l_41 [2317] &  i[1819]);
assign l_40[1160]    = ( l_41 [2318] & !i[1819]) | ( l_41 [2319] &  i[1819]);
assign l_40[1161]    = ( l_41 [2320] & !i[1819]) | ( l_41 [2321] &  i[1819]);
assign l_40[1162]    = ( l_41 [2322] & !i[1819]) | ( l_41 [2323] &  i[1819]);
assign l_40[1163]    = ( l_41 [2324] & !i[1819]) | ( l_41 [2325] &  i[1819]);
assign l_40[1164]    = ( l_41 [2326] & !i[1819]) | ( l_41 [2327] &  i[1819]);
assign l_40[1165]    = ( l_41 [2328] & !i[1819]) | ( l_41 [2329] &  i[1819]);
assign l_40[1166]    = ( l_41 [2330] & !i[1819]) | ( l_41 [2331] &  i[1819]);
assign l_40[1167]    = ( l_41 [2332] & !i[1819]) | ( l_41 [2333] &  i[1819]);
assign l_40[1168]    = ( l_41 [2334] & !i[1819]) | ( l_41 [2335] &  i[1819]);
assign l_40[1169]    = ( l_41 [2336] & !i[1819]) | ( l_41 [2337] &  i[1819]);
assign l_40[1170]    = ( l_41 [2338] & !i[1819]) | ( l_41 [2339] &  i[1819]);
assign l_40[1171]    = ( l_41 [2340] & !i[1819]) | ( l_41 [2341] &  i[1819]);
assign l_40[1172]    = ( l_41 [2342] & !i[1819]) | ( l_41 [2343] &  i[1819]);
assign l_40[1173]    = ( l_41 [2344] & !i[1819]) | ( l_41 [2345] &  i[1819]);
assign l_40[1174]    = ( l_41 [2346] & !i[1819]) | ( l_41 [2347] &  i[1819]);
assign l_40[1175]    = ( l_41 [2348] & !i[1819]) | ( l_41 [2349] &  i[1819]);
assign l_40[1176]    = ( l_41 [2350] & !i[1819]) | ( l_41 [2351] &  i[1819]);
assign l_40[1177]    = ( l_41 [2352] & !i[1819]) | ( l_41 [2353] &  i[1819]);
assign l_40[1178]    = ( l_41 [2354] & !i[1819]) | ( l_41 [2355] &  i[1819]);
assign l_40[1179]    = ( l_41 [2356] & !i[1819]) | ( l_41 [2357] &  i[1819]);
assign l_40[1180]    = ( l_41 [2358] & !i[1819]) | ( l_41 [2359] &  i[1819]);
assign l_40[1181]    = ( l_41 [2360] & !i[1819]) | ( l_41 [2361] &  i[1819]);
assign l_40[1182]    = ( l_41 [2362] & !i[1819]) | ( l_41 [2363] &  i[1819]);
assign l_40[1183]    = ( l_41 [2364] & !i[1819]) | ( l_41 [2365] &  i[1819]);
assign l_40[1184]    = ( l_41 [2366] & !i[1819]) | ( l_41 [2367] &  i[1819]);
assign l_40[1185]    = ( l_41 [2368] & !i[1819]) | ( l_41 [2369] &  i[1819]);
assign l_40[1186]    = ( l_41 [2370] & !i[1819]) | ( l_41 [2371] &  i[1819]);
assign l_40[1187]    = ( l_41 [2372] & !i[1819]) | ( l_41 [2373] &  i[1819]);
assign l_40[1188]    = ( l_41 [2374] & !i[1819]) | ( l_41 [2375] &  i[1819]);
assign l_40[1189]    = ( l_41 [2376] & !i[1819]) | ( l_41 [2377] &  i[1819]);
assign l_40[1190]    = ( l_41 [2378] & !i[1819]) | ( l_41 [2379] &  i[1819]);
assign l_40[1191]    = ( l_41 [2380] & !i[1819]) | ( l_41 [2381] &  i[1819]);
assign l_40[1192]    = ( l_41 [2382] & !i[1819]) | ( l_41 [2383] &  i[1819]);
assign l_40[1193]    = ( l_41 [2384] & !i[1819]) | ( l_41 [2385] &  i[1819]);
assign l_40[1194]    = ( l_41 [2386] & !i[1819]) | ( l_41 [2387] &  i[1819]);
assign l_40[1195]    = ( l_41 [2388] & !i[1819]) | ( l_41 [2389] &  i[1819]);
assign l_40[1196]    = ( l_41 [2390] & !i[1819]) | ( l_41 [2391] &  i[1819]);
assign l_40[1197]    = ( l_41 [2392] & !i[1819]) | ( l_41 [2393] &  i[1819]);
assign l_40[1198]    = ( l_41 [2394] & !i[1819]) | ( l_41 [2395] &  i[1819]);
assign l_40[1199]    = ( l_41 [2396] & !i[1819]) | ( l_41 [2397] &  i[1819]);
assign l_40[1200]    = ( l_41 [2398] & !i[1819]) | ( l_41 [2399] &  i[1819]);
assign l_40[1201]    = ( l_41 [2400] & !i[1819]) | ( l_41 [2401] &  i[1819]);
assign l_40[1202]    = ( l_41 [2402] & !i[1819]) | ( l_41 [2403] &  i[1819]);
assign l_40[1203]    = ( l_41 [2404] & !i[1819]) | ( l_41 [2405] &  i[1819]);
assign l_40[1204]    = ( l_41 [2406] & !i[1819]) | ( l_41 [2407] &  i[1819]);
assign l_40[1205]    = ( l_41 [2408] & !i[1819]) | ( l_41 [2409] &  i[1819]);
assign l_40[1206]    = ( l_41 [2410] & !i[1819]) | ( l_41 [2411] &  i[1819]);
assign l_40[1207]    = ( l_41 [2412] & !i[1819]) | ( l_41 [2413] &  i[1819]);
assign l_40[1208]    = ( l_41 [2414] & !i[1819]) | ( l_41 [2415] &  i[1819]);
assign l_40[1209]    = ( l_41 [2416] & !i[1819]) | ( l_41 [2417] &  i[1819]);
assign l_40[1210]    = ( l_41 [2418] & !i[1819]) | ( l_41 [2419] &  i[1819]);
assign l_40[1211]    = ( l_41 [2420] & !i[1819]) | ( l_41 [2421] &  i[1819]);
assign l_40[1212]    = ( l_41 [2422] & !i[1819]) | ( l_41 [2423] &  i[1819]);
assign l_40[1213]    = ( l_41 [2424] & !i[1819]) | ( l_41 [2425] &  i[1819]);
assign l_40[1214]    = ( l_41 [2426] & !i[1819]) | ( l_41 [2427] &  i[1819]);
assign l_40[1215]    = ( l_41 [2428] & !i[1819]) | ( l_41 [2429] &  i[1819]);
assign l_40[1216]    = ( l_41 [2430] & !i[1819]) | ( l_41 [2431] &  i[1819]);
assign l_40[1217]    = ( l_41 [2432] & !i[1819]) | ( l_41 [2433] &  i[1819]);
assign l_40[1218]    = ( l_41 [2434] & !i[1819]) | ( l_41 [2435] &  i[1819]);
assign l_40[1219]    = ( l_41 [2436] & !i[1819]) | ( l_41 [2437] &  i[1819]);
assign l_40[1220]    = ( l_41 [2438] & !i[1819]) | ( l_41 [2439] &  i[1819]);
assign l_40[1221]    = ( l_41 [2440] & !i[1819]) | ( l_41 [2441] &  i[1819]);
assign l_40[1222]    = ( l_41 [2442] & !i[1819]) | ( l_41 [2443] &  i[1819]);
assign l_40[1223]    = ( l_41 [2444] & !i[1819]) | ( l_41 [2445] &  i[1819]);
assign l_40[1224]    = ( l_41 [2446] & !i[1819]) | ( l_41 [2447] &  i[1819]);
assign l_40[1225]    = ( l_41 [2448] & !i[1819]) | ( l_41 [2449] &  i[1819]);
assign l_40[1226]    = ( l_41 [2450] & !i[1819]) | ( l_41 [2451] &  i[1819]);
assign l_40[1227]    = ( l_41 [2452] & !i[1819]) | ( l_41 [2453] &  i[1819]);
assign l_40[1228]    = ( l_41 [2454] & !i[1819]) | ( l_41 [2455] &  i[1819]);
assign l_40[1229]    = ( l_41 [2456] & !i[1819]) | ( l_41 [2457] &  i[1819]);
assign l_40[1230]    = ( l_41 [2458] & !i[1819]) | ( l_41 [2459] &  i[1819]);
assign l_40[1231]    = ( l_41 [2460] & !i[1819]) | ( l_41 [2461] &  i[1819]);
assign l_40[1232]    = ( l_41 [2462] & !i[1819]) | ( l_41 [2463] &  i[1819]);
assign l_40[1233]    = ( l_41 [2464] & !i[1819]) | ( l_41 [2465] &  i[1819]);
assign l_40[1234]    = ( l_41 [2466] & !i[1819]) | ( l_41 [2467] &  i[1819]);
assign l_40[1235]    = ( l_41 [2468] & !i[1819]) | ( l_41 [2469] &  i[1819]);
assign l_40[1236]    = ( l_41 [2470] & !i[1819]) | ( l_41 [2471] &  i[1819]);
assign l_40[1237]    = ( l_41 [2472] & !i[1819]) | ( l_41 [2473] &  i[1819]);
assign l_40[1238]    = ( l_41 [2474] & !i[1819]) | ( l_41 [2475] &  i[1819]);
assign l_40[1239]    = ( l_41 [2476] & !i[1819]) | ( l_41 [2477] &  i[1819]);
assign l_40[1240]    = ( l_41 [2478] & !i[1819]) | ( l_41 [2479] &  i[1819]);
assign l_40[1241]    = ( l_41 [2480] & !i[1819]) | ( l_41 [2481] &  i[1819]);
assign l_40[1242]    = ( l_41 [2482] & !i[1819]) | ( l_41 [2483] &  i[1819]);
assign l_40[1243]    = ( l_41 [2484] & !i[1819]) | ( l_41 [2485] &  i[1819]);
assign l_40[1244]    = ( l_41 [2486] & !i[1819]) | ( l_41 [2487] &  i[1819]);
assign l_40[1245]    = ( l_41 [2488] & !i[1819]) | ( l_41 [2489] &  i[1819]);
assign l_40[1246]    = ( l_41 [2490] & !i[1819]) | ( l_41 [2491] &  i[1819]);
assign l_40[1247]    = ( l_41 [2492] & !i[1819]) | ( l_41 [2493] &  i[1819]);
assign l_40[1248]    = ( l_41 [2494] & !i[1819]) | ( l_41 [2495] &  i[1819]);
assign l_40[1249]    = ( l_41 [2496] & !i[1819]) | ( l_41 [2497] &  i[1819]);
assign l_40[1250]    = ( l_41 [2498] & !i[1819]) | ( l_41 [2499] &  i[1819]);
assign l_40[1251]    = ( l_41 [2500] & !i[1819]) | ( l_41 [2501] &  i[1819]);
assign l_40[1252]    = ( l_41 [2502] & !i[1819]) | ( l_41 [2503] &  i[1819]);
assign l_40[1253]    = ( l_41 [2504] & !i[1819]) | ( l_41 [2505] &  i[1819]);
assign l_40[1254]    = ( l_41 [2506] & !i[1819]) | ( l_41 [2507] &  i[1819]);
assign l_40[1255]    = ( l_41 [2508] & !i[1819]) | ( l_41 [2509] &  i[1819]);
assign l_40[1256]    = ( l_41 [2510] & !i[1819]) | ( l_41 [2511] &  i[1819]);
assign l_40[1257]    = ( l_41 [2512] & !i[1819]) | ( l_41 [2513] &  i[1819]);
assign l_40[1258]    = ( l_41 [2514] & !i[1819]) | ( l_41 [2515] &  i[1819]);
assign l_40[1259]    = ( l_41 [2516] & !i[1819]) | ( l_41 [2517] &  i[1819]);
assign l_40[1260]    = ( l_41 [2518] & !i[1819]) | ( l_41 [2519] &  i[1819]);
assign l_40[1261]    = ( l_41 [2520] & !i[1819]) | ( l_41 [2521] &  i[1819]);
assign l_40[1262]    = ( l_41 [2522] & !i[1819]) | ( l_41 [2523] &  i[1819]);
assign l_40[1263]    = ( l_41 [2524] & !i[1819]) | ( l_41 [2525] &  i[1819]);
assign l_40[1264]    = ( l_41 [2526] & !i[1819]) | ( l_41 [2527] &  i[1819]);
assign l_40[1265]    = ( l_41 [2528] & !i[1819]) | ( l_41 [2529] &  i[1819]);
assign l_40[1266]    = ( l_41 [2530] & !i[1819]) | ( l_41 [2531] &  i[1819]);
assign l_40[1267]    = ( l_41 [2532] & !i[1819]) | ( l_41 [2533] &  i[1819]);
assign l_40[1268]    = ( l_41 [2534] & !i[1819]) | ( l_41 [2535] &  i[1819]);
assign l_40[1269]    = ( l_41 [2536] & !i[1819]) | ( l_41 [2537] &  i[1819]);
assign l_40[1270]    = ( l_41 [2538] & !i[1819]) | ( l_41 [2539] &  i[1819]);
assign l_40[1271]    = ( l_41 [2540] & !i[1819]) | ( l_41 [2541] &  i[1819]);
assign l_40[1272]    = ( l_41 [2542] & !i[1819]) | ( l_41 [2543] &  i[1819]);
assign l_40[1273]    = ( l_41 [2544] & !i[1819]) | ( l_41 [2545] &  i[1819]);
assign l_40[1274]    = ( l_41 [2546] & !i[1819]) | ( l_41 [2547] &  i[1819]);
assign l_40[1275]    = ( l_41 [2548] & !i[1819]) | ( l_41 [2549] &  i[1819]);
assign l_40[1276]    = ( l_41 [2550] & !i[1819]) | ( l_41 [2551] &  i[1819]);
assign l_40[1277]    = ( l_41 [2552] & !i[1819]) | ( l_41 [2553] &  i[1819]);
assign l_40[1278]    = ( l_41 [2554] & !i[1819]) | ( l_41 [2555] &  i[1819]);
assign l_40[1279]    = ( l_41 [2556] & !i[1819]) | ( l_41 [2557] &  i[1819]);
assign l_40[1280]    = ( l_41 [2558] & !i[1819]) | ( l_41 [2559] &  i[1819]);
assign l_40[1281]    = ( l_41 [2560] & !i[1819]) | ( l_41 [2561] &  i[1819]);
assign l_40[1282]    = ( l_41 [2562] & !i[1819]) | ( l_41 [2563] &  i[1819]);
assign l_40[1283]    = ( l_41 [2564] & !i[1819]) | ( l_41 [2565] &  i[1819]);
assign l_40[1284]    = ( l_41 [2566] & !i[1819]) | ( l_41 [2567] &  i[1819]);
assign l_40[1285]    = ( l_41 [2568] & !i[1819]) | ( l_41 [2569] &  i[1819]);
assign l_40[1286]    = ( l_41 [2570] & !i[1819]) | ( l_41 [2571] &  i[1819]);
assign l_40[1287]    = ( l_41 [2572] & !i[1819]) | ( l_41 [2573] &  i[1819]);
assign l_40[1288]    = ( l_41 [2574] & !i[1819]) | ( l_41 [2575] &  i[1819]);
assign l_40[1289]    = ( l_41 [2576] & !i[1819]) | ( l_41 [2577] &  i[1819]);
assign l_40[1290]    = ( l_41 [2578] & !i[1819]) | ( l_41 [2579] &  i[1819]);
assign l_40[1291]    = ( l_41 [2580] & !i[1819]) | ( l_41 [2581] &  i[1819]);
assign l_40[1292]    = ( l_41 [2582] & !i[1819]) | ( l_41 [2583] &  i[1819]);
assign l_40[1293]    = ( l_41 [2584] & !i[1819]) | ( l_41 [2585] &  i[1819]);
assign l_40[1294]    = ( l_41 [2586] & !i[1819]) | ( l_41 [2587] &  i[1819]);
assign l_40[1295]    = ( l_41 [2588] & !i[1819]) | ( l_41 [2589] &  i[1819]);
assign l_40[1296]    = ( l_41 [2590] & !i[1819]) | ( l_41 [2591] &  i[1819]);
assign l_40[1297]    = ( l_41 [2592] & !i[1819]) | ( l_41 [2593] &  i[1819]);
assign l_40[1298]    = ( l_41 [2594] & !i[1819]) | ( l_41 [2595] &  i[1819]);
assign l_40[1299]    = ( l_41 [2596] & !i[1819]) | ( l_41 [2597] &  i[1819]);
assign l_40[1300]    = ( l_41 [2598] & !i[1819]) | ( l_41 [2599] &  i[1819]);
assign l_40[1301]    = ( l_41 [2600] & !i[1819]) | ( l_41 [2601] &  i[1819]);
assign l_40[1302]    = ( l_41 [2602] & !i[1819]) | ( l_41 [2603] &  i[1819]);
assign l_40[1303]    = ( l_41 [2604] & !i[1819]) | ( l_41 [2605] &  i[1819]);
assign l_40[1304]    = ( l_41 [2606] & !i[1819]) | ( l_41 [2607] &  i[1819]);
assign l_40[1305]    = ( l_41 [2608] & !i[1819]) | ( l_41 [2609] &  i[1819]);
assign l_40[1306]    = ( l_41 [2610] & !i[1819]) | ( l_41 [2611] &  i[1819]);
assign l_40[1307]    = ( l_41 [2612] & !i[1819]) | ( l_41 [2613] &  i[1819]);
assign l_40[1308]    = ( l_41 [2614] & !i[1819]) | ( l_41 [2615] &  i[1819]);
assign l_40[1309]    = ( l_41 [2616] & !i[1819]) | ( l_41 [2617] &  i[1819]);
assign l_40[1310]    = ( l_41 [2618] & !i[1819]) | ( l_41 [2619] &  i[1819]);
assign l_40[1311]    = ( l_41 [2620] & !i[1819]) | ( l_41 [2621] &  i[1819]);
assign l_40[1312]    = ( l_41 [2622] & !i[1819]) | ( l_41 [2623] &  i[1819]);
assign l_40[1313]    = ( l_41 [2624] & !i[1819]) | ( l_41 [2625] &  i[1819]);
assign l_40[1314]    = ( l_41 [2626] & !i[1819]) | ( l_41 [2627] &  i[1819]);
assign l_40[1315]    = ( l_41 [2628] & !i[1819]) | ( l_41 [2629] &  i[1819]);
assign l_40[1316]    = ( l_41 [2630] & !i[1819]) | ( l_41 [2631] &  i[1819]);
assign l_40[1317]    = ( l_41 [2632] & !i[1819]) | ( l_41 [2633] &  i[1819]);
assign l_40[1318]    = ( l_41 [2634] & !i[1819]) | ( l_41 [2635] &  i[1819]);
assign l_40[1319]    = ( l_41 [2636] & !i[1819]) | ( l_41 [2637] &  i[1819]);
assign l_40[1320]    = ( l_41 [2638] & !i[1819]) | ( l_41 [2639] &  i[1819]);
assign l_40[1321]    = ( l_41 [2640] & !i[1819]) | ( l_41 [2641] &  i[1819]);
assign l_40[1322]    = ( l_41 [2642] & !i[1819]) | ( l_41 [2643] &  i[1819]);
assign l_40[1323]    = ( l_41 [2644] & !i[1819]) | ( l_41 [2645] &  i[1819]);
assign l_40[1324]    = ( l_41 [2646] & !i[1819]) | ( l_41 [2647] &  i[1819]);
assign l_40[1325]    = ( l_41 [2648] & !i[1819]) | ( l_41 [2649] &  i[1819]);
assign l_40[1326]    = ( l_41 [2650] & !i[1819]) | ( l_41 [2651] &  i[1819]);
assign l_40[1327]    = ( l_41 [2652] & !i[1819]) | ( l_41 [2653] &  i[1819]);
assign l_40[1328]    = ( l_41 [2654] & !i[1819]) | ( l_41 [2655] &  i[1819]);
assign l_40[1329]    = ( l_41 [2656] & !i[1819]) | ( l_41 [2657] &  i[1819]);
assign l_40[1330]    = ( l_41 [2658] & !i[1819]) | ( l_41 [2659] &  i[1819]);
assign l_40[1331]    = ( l_41 [2660] & !i[1819]) | ( l_41 [2661] &  i[1819]);
assign l_40[1332]    = ( l_41 [2662] & !i[1819]) | ( l_41 [2663] &  i[1819]);
assign l_40[1333]    = ( l_41 [2664] & !i[1819]) | ( l_41 [2665] &  i[1819]);
assign l_40[1334]    = ( l_41 [2666] & !i[1819]) | ( l_41 [2667] &  i[1819]);
assign l_40[1335]    = ( l_41 [2668] & !i[1819]) | ( l_41 [2669] &  i[1819]);
assign l_40[1336]    = ( l_41 [2670] & !i[1819]) | ( l_41 [2671] &  i[1819]);
assign l_40[1337]    = ( l_41 [2672] & !i[1819]) | ( l_41 [2673] &  i[1819]);
assign l_40[1338]    = ( l_41 [2674] & !i[1819]) | ( l_41 [2675] &  i[1819]);
assign l_40[1339]    = ( l_41 [2676] & !i[1819]) | ( l_41 [2677] &  i[1819]);
assign l_40[1340]    = ( l_41 [2678] & !i[1819]) | ( l_41 [2679] &  i[1819]);
assign l_40[1341]    = ( l_41 [2680] & !i[1819]) | ( l_41 [2681] &  i[1819]);
assign l_40[1342]    = ( l_41 [2682] & !i[1819]) | ( l_41 [2683] &  i[1819]);
assign l_40[1343]    = ( l_41 [2684] & !i[1819]) | ( l_41 [2685] &  i[1819]);
assign l_40[1344]    = ( l_41 [2686] & !i[1819]) | ( l_41 [2687] &  i[1819]);
assign l_40[1345]    = ( l_41 [2688] & !i[1819]) | ( l_41 [2689] &  i[1819]);
assign l_40[1346]    = ( l_41 [2690] & !i[1819]) | ( l_41 [2691] &  i[1819]);
assign l_40[1347]    = ( l_41 [2692] & !i[1819]) | ( l_41 [2693] &  i[1819]);
assign l_40[1348]    = ( l_41 [2694] & !i[1819]) | ( l_41 [2695] &  i[1819]);
assign l_40[1349]    = ( l_41 [2696] & !i[1819]) | ( l_41 [2697] &  i[1819]);
assign l_40[1350]    = ( l_41 [2698] & !i[1819]) | ( l_41 [2699] &  i[1819]);
assign l_40[1351]    = ( l_41 [2700] & !i[1819]) | ( l_41 [2701] &  i[1819]);
assign l_40[1352]    = ( l_41 [2702] & !i[1819]) | ( l_41 [2703] &  i[1819]);
assign l_40[1353]    = ( l_41 [2704] & !i[1819]) | ( l_41 [2705] &  i[1819]);
assign l_40[1354]    = ( l_41 [2706] & !i[1819]) | ( l_41 [2707] &  i[1819]);
assign l_40[1355]    = ( l_41 [2708] & !i[1819]) | ( l_41 [2709] &  i[1819]);
assign l_40[1356]    = ( l_41 [2710] & !i[1819]) | ( l_41 [2711] &  i[1819]);
assign l_40[1357]    = ( l_41 [2712] & !i[1819]) | ( l_41 [2713] &  i[1819]);
assign l_40[1358]    = ( l_41 [2714] & !i[1819]) | ( l_41 [2715] &  i[1819]);
assign l_40[1359]    = ( l_41 [2716] & !i[1819]) | ( l_41 [2717] &  i[1819]);
assign l_40[1360]    = ( l_41 [2718] & !i[1819]) | ( l_41 [2719] &  i[1819]);
assign l_40[1361]    = ( l_41 [2720] & !i[1819]) | ( l_41 [2721] &  i[1819]);
assign l_40[1362]    = ( l_41 [2722] & !i[1819]) | ( l_41 [2723] &  i[1819]);
assign l_40[1363]    = ( l_41 [2724] & !i[1819]) | ( l_41 [2725] &  i[1819]);
assign l_40[1364]    = ( l_41 [2726] & !i[1819]) | ( l_41 [2727] &  i[1819]);
assign l_40[1365]    = ( l_41 [2728] & !i[1819]) | ( l_41 [2729] &  i[1819]);
assign l_40[1366]    = ( l_41 [2730] & !i[1819]) | ( l_41 [2731] &  i[1819]);
assign l_40[1367]    = ( l_41 [2732] & !i[1819]) | ( l_41 [2733] &  i[1819]);
assign l_40[1368]    = ( l_41 [2734] & !i[1819]) | ( l_41 [2735] &  i[1819]);
assign l_40[1369]    = ( l_41 [2736] & !i[1819]) | ( l_41 [2737] &  i[1819]);
assign l_40[1370]    = ( l_41 [2738] & !i[1819]) | ( l_41 [2739] &  i[1819]);
assign l_40[1371]    = ( l_41 [2740] & !i[1819]) | ( l_41 [2741] &  i[1819]);
assign l_40[1372]    = ( l_41 [2742] & !i[1819]) | ( l_41 [2743] &  i[1819]);
assign l_40[1373]    = ( l_41 [2744] & !i[1819]) | ( l_41 [2745] &  i[1819]);
assign l_40[1374]    = ( l_41 [2746] & !i[1819]) | ( l_41 [2747] &  i[1819]);
assign l_40[1375]    = ( l_41 [2748] & !i[1819]) | ( l_41 [2749] &  i[1819]);
assign l_40[1376]    = ( l_41 [2750] & !i[1819]) | ( l_41 [2751] &  i[1819]);
assign l_40[1377]    = ( l_41 [2752] & !i[1819]) | ( l_41 [2753] &  i[1819]);
assign l_40[1378]    = ( l_41 [2754] & !i[1819]) | ( l_41 [2755] &  i[1819]);
assign l_40[1379]    = ( l_41 [2756] & !i[1819]) | ( l_41 [2757] &  i[1819]);
assign l_40[1380]    = ( l_41 [2758] & !i[1819]) | ( l_41 [2759] &  i[1819]);
assign l_40[1381]    = ( l_41 [2760] & !i[1819]) | ( l_41 [2761] &  i[1819]);
assign l_40[1382]    = ( l_41 [2762] & !i[1819]) | ( l_41 [2763] &  i[1819]);
assign l_40[1383]    = ( l_41 [2764] & !i[1819]) | ( l_41 [2765] &  i[1819]);
assign l_40[1384]    = ( l_41 [2766] & !i[1819]) | ( l_41 [2767] &  i[1819]);
assign l_40[1385]    = ( l_41 [2768] & !i[1819]) | ( l_41 [2769] &  i[1819]);
assign l_40[1386]    = ( l_41 [2770] & !i[1819]) | ( l_41 [2771] &  i[1819]);
assign l_40[1387]    = ( l_41 [2772] & !i[1819]) | ( l_41 [2773] &  i[1819]);
assign l_40[1388]    = ( l_41 [2774] & !i[1819]) | ( l_41 [2775] &  i[1819]);
assign l_40[1389]    = ( l_41 [2776] & !i[1819]) | ( l_41 [2777] &  i[1819]);
assign l_40[1390]    = ( l_41 [2778] & !i[1819]) | ( l_41 [2779] &  i[1819]);
assign l_40[1391]    = ( l_41 [2780] & !i[1819]) | ( l_41 [2781] &  i[1819]);
assign l_40[1392]    = ( l_41 [2782] & !i[1819]) | ( l_41 [2783] &  i[1819]);
assign l_40[1393]    = ( l_41 [2784] & !i[1819]) | ( l_41 [2785] &  i[1819]);
assign l_40[1394]    = ( l_41 [2786] & !i[1819]) | ( l_41 [2787] &  i[1819]);
assign l_40[1395]    = ( l_41 [2788] & !i[1819]) | ( l_41 [2789] &  i[1819]);
assign l_40[1396]    = ( l_41 [2790] & !i[1819]) | ( l_41 [2791] &  i[1819]);
assign l_40[1397]    = ( l_41 [2792] & !i[1819]) | ( l_41 [2793] &  i[1819]);
assign l_40[1398]    = ( l_41 [2794] & !i[1819]) | ( l_41 [2795] &  i[1819]);
assign l_40[1399]    = ( l_41 [2796] & !i[1819]) | ( l_41 [2797] &  i[1819]);
assign l_40[1400]    = ( l_41 [2798] & !i[1819]) | ( l_41 [2799] &  i[1819]);
assign l_40[1401]    = ( l_41 [2800] & !i[1819]) | ( l_41 [2801] &  i[1819]);
assign l_40[1402]    = ( l_41 [2802] & !i[1819]) | ( l_41 [2803] &  i[1819]);
assign l_40[1403]    = ( l_41 [2804] & !i[1819]) | ( l_41 [2805] &  i[1819]);
assign l_40[1404]    = ( l_41 [2806] & !i[1819]) | ( l_41 [2807] &  i[1819]);
assign l_40[1405]    = ( l_41 [2808] & !i[1819]) | ( l_41 [2809] &  i[1819]);
assign l_40[1406]    = ( l_41 [2810] & !i[1819]) | ( l_41 [2811] &  i[1819]);
assign l_40[1407]    = ( l_41 [2812] & !i[1819]) | ( l_41 [2813] &  i[1819]);
assign l_40[1408]    = ( l_41 [2814] & !i[1819]) | ( l_41 [2815] &  i[1819]);
assign l_40[1409]    = ( l_41 [2816] & !i[1819]) | ( l_41 [2817] &  i[1819]);
assign l_40[1410]    = ( l_41 [2818] & !i[1819]) | ( l_41 [2819] &  i[1819]);
assign l_40[1411]    = ( l_41 [2820] & !i[1819]) | ( l_41 [2821] &  i[1819]);
assign l_40[1412]    = ( l_41 [2822] & !i[1819]) | ( l_41 [2823] &  i[1819]);
assign l_40[1413]    = ( l_41 [2824] & !i[1819]) | ( l_41 [2825] &  i[1819]);
assign l_40[1414]    = ( l_41 [2826] & !i[1819]) | ( l_41 [2827] &  i[1819]);
assign l_40[1415]    = ( l_41 [2828] & !i[1819]) | ( l_41 [2829] &  i[1819]);
assign l_40[1416]    = ( l_41 [2830] & !i[1819]) | ( l_41 [2831] &  i[1819]);
assign l_40[1417]    = ( l_41 [2832] & !i[1819]) | ( l_41 [2833] &  i[1819]);
assign l_40[1418]    = ( l_41 [2834] & !i[1819]) | ( l_41 [2835] &  i[1819]);
assign l_40[1419]    = ( l_41 [2836] & !i[1819]) | ( l_41 [2837] &  i[1819]);
assign l_40[1420]    = ( l_41 [2838] & !i[1819]) | ( l_41 [2839] &  i[1819]);
assign l_40[1421]    = ( l_41 [2840] & !i[1819]) | ( l_41 [2841] &  i[1819]);
assign l_40[1422]    = ( l_41 [2842] & !i[1819]) | ( l_41 [2843] &  i[1819]);
assign l_40[1423]    = ( l_41 [2844] & !i[1819]) | ( l_41 [2845] &  i[1819]);
assign l_40[1424]    = ( l_41 [2846] & !i[1819]) | ( l_41 [2847] &  i[1819]);
assign l_40[1425]    = ( l_41 [2848] & !i[1819]) | ( l_41 [2849] &  i[1819]);
assign l_40[1426]    = ( l_41 [2850] & !i[1819]) | ( l_41 [2851] &  i[1819]);
assign l_40[1427]    = ( l_41 [2852] & !i[1819]) | ( l_41 [2853] &  i[1819]);
assign l_40[1428]    = ( l_41 [2854] & !i[1819]) | ( l_41 [2855] &  i[1819]);
assign l_40[1429]    = ( l_41 [2856] & !i[1819]) | ( l_41 [2857] &  i[1819]);
assign l_40[1430]    = ( l_41 [2858] & !i[1819]) | ( l_41 [2859] &  i[1819]);
assign l_40[1431]    = ( l_41 [2860] & !i[1819]) | ( l_41 [2861] &  i[1819]);
assign l_40[1432]    = ( l_41 [2862] & !i[1819]) | ( l_41 [2863] &  i[1819]);
assign l_40[1433]    = ( l_41 [2864] & !i[1819]) | ( l_41 [2865] &  i[1819]);
assign l_40[1434]    = ( l_41 [2866] & !i[1819]) | ( l_41 [2867] &  i[1819]);
assign l_40[1435]    = ( l_41 [2868] & !i[1819]) | ( l_41 [2869] &  i[1819]);
assign l_40[1436]    = ( l_41 [2870] & !i[1819]) | ( l_41 [2871] &  i[1819]);
assign l_40[1437]    = ( l_41 [2872] & !i[1819]) | ( l_41 [2873] &  i[1819]);
assign l_40[1438]    = ( l_41 [2874] & !i[1819]) | ( l_41 [2875] &  i[1819]);
assign l_40[1439]    = ( l_41 [2876] & !i[1819]) | ( l_41 [2877] &  i[1819]);
assign l_40[1440]    = ( l_41 [2878] & !i[1819]) | ( l_41 [2879] &  i[1819]);
assign l_40[1441]    = ( l_41 [2880] & !i[1819]) | ( l_41 [2881] &  i[1819]);
assign l_40[1442]    = ( l_41 [2882] & !i[1819]) | ( l_41 [2883] &  i[1819]);
assign l_40[1443]    = ( l_41 [2884] & !i[1819]) | ( l_41 [2885] &  i[1819]);
assign l_40[1444]    = ( l_41 [2886] & !i[1819]) | ( l_41 [2887] &  i[1819]);
assign l_40[1445]    = ( l_41 [2888] & !i[1819]) | ( l_41 [2889] &  i[1819]);
assign l_40[1446]    = ( l_41 [2890] & !i[1819]) | ( l_41 [2891] &  i[1819]);
assign l_40[1447]    = ( l_41 [2892] & !i[1819]) | ( l_41 [2893] &  i[1819]);
assign l_40[1448]    = ( l_41 [2894] & !i[1819]) | ( l_41 [2895] &  i[1819]);
assign l_40[1449]    = ( l_41 [2896] & !i[1819]) | ( l_41 [2897] &  i[1819]);
assign l_40[1450]    = ( l_41 [2898] & !i[1819]) | ( l_41 [2899] &  i[1819]);
assign l_40[1451]    = ( l_41 [2900] & !i[1819]) | ( l_41 [2901] &  i[1819]);
assign l_40[1452]    = ( l_41 [2902] & !i[1819]) | ( l_41 [2903] &  i[1819]);
assign l_40[1453]    = ( l_41 [2904] & !i[1819]) | ( l_41 [2905] &  i[1819]);
assign l_40[1454]    = ( l_41 [2906] & !i[1819]) | ( l_41 [2907] &  i[1819]);
assign l_40[1455]    = ( l_41 [2908] & !i[1819]) | ( l_41 [2909] &  i[1819]);
assign l_40[1456]    = ( l_41 [2910] & !i[1819]) | ( l_41 [2911] &  i[1819]);
assign l_40[1457]    = ( l_41 [2912] & !i[1819]) | ( l_41 [2913] &  i[1819]);
assign l_40[1458]    = ( l_41 [2914] & !i[1819]) | ( l_41 [2915] &  i[1819]);
assign l_40[1459]    = ( l_41 [2916] & !i[1819]) | ( l_41 [2917] &  i[1819]);
assign l_40[1460]    = ( l_41 [2918] & !i[1819]) | ( l_41 [2919] &  i[1819]);
assign l_40[1461]    = ( l_41 [2920] & !i[1819]) | ( l_41 [2921] &  i[1819]);
assign l_40[1462]    = ( l_41 [2922] & !i[1819]) | ( l_41 [2923] &  i[1819]);
assign l_40[1463]    = ( l_41 [2924] & !i[1819]) | ( l_41 [2925] &  i[1819]);
assign l_40[1464]    = ( l_41 [2926] & !i[1819]) | ( l_41 [2927] &  i[1819]);
assign l_40[1465]    = ( l_41 [2928] & !i[1819]) | ( l_41 [2929] &  i[1819]);
assign l_40[1466]    = ( l_41 [2930] & !i[1819]) | ( l_41 [2931] &  i[1819]);
assign l_40[1467]    = ( l_41 [2932] & !i[1819]) | ( l_41 [2933] &  i[1819]);
assign l_40[1468]    = ( l_41 [2934] & !i[1819]) | ( l_41 [2935] &  i[1819]);
assign l_40[1469]    = ( l_41 [2936] & !i[1819]) | ( l_41 [2937] &  i[1819]);
assign l_40[1470]    = ( l_41 [2938] & !i[1819]) | ( l_41 [2939] &  i[1819]);
assign l_40[1471]    = ( l_41 [2940] & !i[1819]) | ( l_41 [2941] &  i[1819]);
assign l_40[1472]    = ( l_41 [2942] & !i[1819]) | ( l_41 [2943] &  i[1819]);
assign l_40[1473]    = ( l_41 [2944] & !i[1819]) | ( l_41 [2945] &  i[1819]);
assign l_40[1474]    = ( l_41 [2946] & !i[1819]) | ( l_41 [2947] &  i[1819]);
assign l_40[1475]    = ( l_41 [2948] & !i[1819]) | ( l_41 [2949] &  i[1819]);
assign l_40[1476]    = ( l_41 [2950] & !i[1819]) | ( l_41 [2951] &  i[1819]);
assign l_40[1477]    = ( l_41 [2952] & !i[1819]) | ( l_41 [2953] &  i[1819]);
assign l_40[1478]    = ( l_41 [2954] & !i[1819]) | ( l_41 [2955] &  i[1819]);
assign l_40[1479]    = ( l_41 [2956] & !i[1819]) | ( l_41 [2957] &  i[1819]);
assign l_40[1480]    = ( l_41 [2958] & !i[1819]) | ( l_41 [2959] &  i[1819]);
assign l_40[1481]    = ( l_41 [2960] & !i[1819]) | ( l_41 [2961] &  i[1819]);
assign l_40[1482]    = ( l_41 [2962] & !i[1819]) | ( l_41 [2963] &  i[1819]);
assign l_40[1483]    = ( l_41 [2964] & !i[1819]) | ( l_41 [2965] &  i[1819]);
assign l_40[1484]    = ( l_41 [2966] & !i[1819]) | ( l_41 [2967] &  i[1819]);
assign l_40[1485]    = ( l_41 [2968] & !i[1819]) | ( l_41 [2969] &  i[1819]);
assign l_40[1486]    = ( l_41 [2970] & !i[1819]) | ( l_41 [2971] &  i[1819]);
assign l_40[1487]    = ( l_41 [2972] & !i[1819]) | ( l_41 [2973] &  i[1819]);
assign l_40[1488]    = ( l_41 [2974] & !i[1819]) | ( l_41 [2975] &  i[1819]);
assign l_40[1489]    = ( l_41 [2976] & !i[1819]) | ( l_41 [2977] &  i[1819]);
assign l_40[1490]    = ( l_41 [2978] & !i[1819]) | ( l_41 [2979] &  i[1819]);
assign l_40[1491]    = ( l_41 [2980] & !i[1819]) | ( l_41 [2981] &  i[1819]);
assign l_40[1492]    = ( l_41 [2982] & !i[1819]) | ( l_41 [2983] &  i[1819]);
assign l_40[1493]    = ( l_41 [2984] & !i[1819]) | ( l_41 [2985] &  i[1819]);
assign l_40[1494]    = ( l_41 [2986] & !i[1819]) | ( l_41 [2987] &  i[1819]);
assign l_40[1495]    = ( l_41 [2988] & !i[1819]) | ( l_41 [2989] &  i[1819]);
assign l_40[1496]    = ( l_41 [2990] & !i[1819]) | ( l_41 [2991] &  i[1819]);
assign l_40[1497]    = ( l_41 [2992] & !i[1819]) | ( l_41 [2993] &  i[1819]);
assign l_40[1498]    = ( l_41 [2994] & !i[1819]) | ( l_41 [2995] &  i[1819]);
assign l_40[1499]    = ( l_41 [2996] & !i[1819]) | ( l_41 [2997] &  i[1819]);
assign l_40[1500]    = ( l_41 [2998] & !i[1819]) | ( l_41 [2999] &  i[1819]);
assign l_40[1501]    = ( l_41 [3000] & !i[1819]) | ( l_41 [3001] &  i[1819]);
assign l_40[1502]    = ( l_41 [3002] & !i[1819]) | ( l_41 [3003] &  i[1819]);
assign l_40[1503]    = ( l_41 [3004] & !i[1819]) | ( l_41 [3005] &  i[1819]);
assign l_40[1504]    = ( l_41 [3006] & !i[1819]) | ( l_41 [3007] &  i[1819]);
assign l_40[1505]    = ( l_41 [3008] & !i[1819]) | ( l_41 [3009] &  i[1819]);
assign l_40[1506]    = ( l_41 [3010] & !i[1819]) | ( l_41 [3011] &  i[1819]);
assign l_40[1507]    = ( l_41 [3012] & !i[1819]) | ( l_41 [3013] &  i[1819]);
assign l_40[1508]    = ( l_41 [3014] & !i[1819]) | ( l_41 [3015] &  i[1819]);
assign l_40[1509]    = ( l_41 [3016] & !i[1819]) | ( l_41 [3017] &  i[1819]);
assign l_40[1510]    = ( l_41 [3018] & !i[1819]) | ( l_41 [3019] &  i[1819]);
assign l_40[1511]    = ( l_41 [3020] & !i[1819]) | ( l_41 [3021] &  i[1819]);
assign l_40[1512]    = ( l_41 [3022] & !i[1819]) | ( l_41 [3023] &  i[1819]);
assign l_40[1513]    = ( l_41 [3024] & !i[1819]) | ( l_41 [3025] &  i[1819]);
assign l_40[1514]    = ( l_41 [3026] & !i[1819]) | ( l_41 [3027] &  i[1819]);
assign l_40[1515]    = ( l_41 [3028] & !i[1819]) | ( l_41 [3029] &  i[1819]);
assign l_40[1516]    = ( l_41 [3030] & !i[1819]) | ( l_41 [3031] &  i[1819]);
assign l_40[1517]    = ( l_41 [3032] & !i[1819]) | ( l_41 [3033] &  i[1819]);
assign l_40[1518]    = ( l_41 [3034] & !i[1819]) | ( l_41 [3035] &  i[1819]);
assign l_40[1519]    = ( l_41 [3036] & !i[1819]) | ( l_41 [3037] &  i[1819]);
assign l_40[1520]    = ( l_41 [3038] & !i[1819]) | ( l_41 [3039] &  i[1819]);
assign l_40[1521]    = ( l_41 [3040] & !i[1819]) | ( l_41 [3041] &  i[1819]);
assign l_40[1522]    = ( l_41 [3042] & !i[1819]) | ( l_41 [3043] &  i[1819]);
assign l_40[1523]    = ( l_41 [3044] & !i[1819]) | ( l_41 [3045] &  i[1819]);
assign l_40[1524]    = ( l_41 [3046] & !i[1819]) | ( l_41 [3047] &  i[1819]);
assign l_40[1525]    = ( l_41 [3048] & !i[1819]) | ( l_41 [3049] &  i[1819]);
assign l_40[1526]    = ( l_41 [3050] & !i[1819]) | ( l_41 [3051] &  i[1819]);
assign l_40[1527]    = ( l_41 [3052] & !i[1819]) | ( l_41 [3053] &  i[1819]);
assign l_40[1528]    = ( l_41 [3054] & !i[1819]) | ( l_41 [3055] &  i[1819]);
assign l_40[1529]    = ( l_41 [3056] & !i[1819]) | ( l_41 [3057] &  i[1819]);
assign l_40[1530]    = ( l_41 [3058] & !i[1819]) | ( l_41 [3059] &  i[1819]);
assign l_40[1531]    = ( l_41 [3060] & !i[1819]) | ( l_41 [3061] &  i[1819]);
assign l_40[1532]    = ( l_41 [3062] & !i[1819]) | ( l_41 [3063] &  i[1819]);
assign l_40[1533]    = ( l_41 [3064] & !i[1819]) | ( l_41 [3065] &  i[1819]);
assign l_40[1534]    = ( l_41 [3066] & !i[1819]) | ( l_41 [3067] &  i[1819]);
assign l_40[1535]    = ( l_41 [3068] & !i[1819]) | ( l_41 [3069] &  i[1819]);
assign l_40[1536]    = ( l_41 [3070] & !i[1819]) | ( l_41 [3071] &  i[1819]);
assign l_40[1537]    = ( l_41 [3072] & !i[1819]) | ( l_41 [3073] &  i[1819]);
assign l_40[1538]    = ( l_41 [3074] & !i[1819]) | ( l_41 [3075] &  i[1819]);
assign l_40[1539]    = ( l_41 [3076] & !i[1819]) | ( l_41 [3077] &  i[1819]);
assign l_40[1540]    = ( l_41 [3078] & !i[1819]) | ( l_41 [3079] &  i[1819]);
assign l_40[1541]    = ( l_41 [3080] & !i[1819]) | ( l_41 [3081] &  i[1819]);
assign l_40[1542]    = ( l_41 [3082] & !i[1819]) | ( l_41 [3083] &  i[1819]);
assign l_40[1543]    = ( l_41 [3084] & !i[1819]) | ( l_41 [3085] &  i[1819]);
assign l_40[1544]    = ( l_41 [3086] & !i[1819]) | ( l_41 [3087] &  i[1819]);
assign l_40[1545]    = ( l_41 [3088] & !i[1819]) | ( l_41 [3089] &  i[1819]);
assign l_40[1546]    = ( l_41 [3090] & !i[1819]) | ( l_41 [3091] &  i[1819]);
assign l_40[1547]    = ( l_41 [3092] & !i[1819]) | ( l_41 [3093] &  i[1819]);
assign l_40[1548]    = ( l_41 [3094] & !i[1819]) | ( l_41 [3095] &  i[1819]);
assign l_40[1549]    = ( l_41 [3096] & !i[1819]) | ( l_41 [3097] &  i[1819]);
assign l_40[1550]    = ( l_41 [3098] & !i[1819]) | ( l_41 [3099] &  i[1819]);
assign l_40[1551]    = ( l_41 [3100] & !i[1819]) | ( l_41 [3101] &  i[1819]);
assign l_40[1552]    = ( l_41 [3102] & !i[1819]) | ( l_41 [3103] &  i[1819]);
assign l_40[1553]    = ( l_41 [3104] & !i[1819]) | ( l_41 [3105] &  i[1819]);
assign l_40[1554]    = ( l_41 [3106] & !i[1819]) | ( l_41 [3107] &  i[1819]);
assign l_40[1555]    = ( l_41 [3108] & !i[1819]) | ( l_41 [3109] &  i[1819]);
assign l_40[1556]    = ( l_41 [3110] & !i[1819]) | ( l_41 [3111] &  i[1819]);
assign l_40[1557]    = ( l_41 [3112] & !i[1819]) | ( l_41 [3113] &  i[1819]);
assign l_40[1558]    = ( l_41 [3114] & !i[1819]) | ( l_41 [3115] &  i[1819]);
assign l_40[1559]    = ( l_41 [3116] & !i[1819]) | ( l_41 [3117] &  i[1819]);
assign l_40[1560]    = ( l_41 [3118] & !i[1819]) | ( l_41 [3119] &  i[1819]);
assign l_40[1561]    = ( l_41 [3120] & !i[1819]) | ( l_41 [3121] &  i[1819]);
assign l_40[1562]    = ( l_41 [3122] & !i[1819]) | ( l_41 [3123] &  i[1819]);
assign l_40[1563]    = ( l_41 [3124] & !i[1819]) | ( l_41 [3125] &  i[1819]);
assign l_40[1564]    = ( l_41 [3126] & !i[1819]) | ( l_41 [3127] &  i[1819]);
assign l_40[1565]    = ( l_41 [3128] & !i[1819]) | ( l_41 [3129] &  i[1819]);
assign l_40[1566]    = ( l_41 [3130] & !i[1819]) | ( l_41 [3131] &  i[1819]);
assign l_40[1567]    = ( l_41 [3132] & !i[1819]) | ( l_41 [3133] &  i[1819]);
assign l_40[1568]    = ( l_41 [3134] & !i[1819]) | ( l_41 [3135] &  i[1819]);
assign l_40[1569]    = ( l_41 [3136] & !i[1819]) | ( l_41 [3137] &  i[1819]);
assign l_40[1570]    = ( l_41 [3138] & !i[1819]) | ( l_41 [3139] &  i[1819]);
assign l_40[1571]    = ( l_41 [3140] & !i[1819]) | ( l_41 [3141] &  i[1819]);
assign l_40[1572]    = ( l_41 [3142] & !i[1819]) | ( l_41 [3143] &  i[1819]);
assign l_40[1573]    = ( l_41 [3144] & !i[1819]) | ( l_41 [3145] &  i[1819]);
assign l_40[1574]    = ( l_41 [3146] & !i[1819]) | ( l_41 [3147] &  i[1819]);
assign l_40[1575]    = ( l_41 [3148] & !i[1819]) | ( l_41 [3149] &  i[1819]);
assign l_40[1576]    = ( l_41 [3150] & !i[1819]) | ( l_41 [3151] &  i[1819]);
assign l_40[1577]    = ( l_41 [3152] & !i[1819]) | ( l_41 [3153] &  i[1819]);
assign l_40[1578]    = ( l_41 [3154] & !i[1819]) | ( l_41 [3155] &  i[1819]);
assign l_40[1579]    = ( l_41 [3156] & !i[1819]) | ( l_41 [3157] &  i[1819]);
assign l_40[1580]    = ( l_41 [3158] & !i[1819]) | ( l_41 [3159] &  i[1819]);
assign l_40[1581]    = ( l_41 [3160] & !i[1819]) | ( l_41 [3161] &  i[1819]);
assign l_40[1582]    = ( l_41 [3162] & !i[1819]) | ( l_41 [3163] &  i[1819]);
assign l_40[1583]    = ( l_41 [3164] & !i[1819]) | ( l_41 [3165] &  i[1819]);
assign l_40[1584]    = ( l_41 [3166] & !i[1819]) | ( l_41 [3167] &  i[1819]);
assign l_40[1585]    = ( l_41 [3168] & !i[1819]) | ( l_41 [3169] &  i[1819]);
assign l_40[1586]    = ( l_41 [3170] & !i[1819]) | ( l_41 [3171] &  i[1819]);
assign l_40[1587]    = ( l_41 [3172] & !i[1819]) | ( l_41 [3173] &  i[1819]);
assign l_40[1588]    = ( l_41 [3174] & !i[1819]) | ( l_41 [3175] &  i[1819]);
assign l_40[1589]    = ( l_41 [3176] & !i[1819]) | ( l_41 [3177] &  i[1819]);
assign l_40[1590]    = ( l_41 [3178] & !i[1819]) | ( l_41 [3179] &  i[1819]);
assign l_40[1591]    = ( l_41 [3180] & !i[1819]) | ( l_41 [3181] &  i[1819]);
assign l_40[1592]    = ( l_41 [3182] & !i[1819]) | ( l_41 [3183] &  i[1819]);
assign l_40[1593]    = ( l_41 [3184] & !i[1819]) | ( l_41 [3185] &  i[1819]);
assign l_40[1594]    = ( l_41 [3186] & !i[1819]) | ( l_41 [3187] &  i[1819]);
assign l_40[1595]    = ( l_41 [3188] & !i[1819]) | ( l_41 [3189] &  i[1819]);
assign l_40[1596]    = ( l_41 [3190] & !i[1819]) | ( l_41 [3191] &  i[1819]);
assign l_40[1597]    = ( l_41 [3192] & !i[1819]) | ( l_41 [3193] &  i[1819]);
assign l_40[1598]    = ( l_41 [3194] & !i[1819]) | ( l_41 [3195] &  i[1819]);
assign l_40[1599]    = ( l_41 [3196] & !i[1819]) | ( l_41 [3197] &  i[1819]);
assign l_40[1600]    = ( l_41 [3198] & !i[1819]) | ( l_41 [3199] &  i[1819]);
assign l_40[1601]    = ( l_41 [3200] & !i[1819]) | ( l_41 [3201] &  i[1819]);
assign l_40[1602]    = ( l_41 [3202] & !i[1819]) | ( l_41 [3203] &  i[1819]);
assign l_40[1603]    = ( l_41 [3204] & !i[1819]) | ( l_41 [3205] &  i[1819]);
assign l_40[1604]    = ( l_41 [3206] & !i[1819]) | ( l_41 [3207] &  i[1819]);
assign l_40[1605]    = ( l_41 [3208] & !i[1819]) | ( l_41 [3209] &  i[1819]);
assign l_40[1606]    = ( l_41 [3210] & !i[1819]) | ( l_41 [3211] &  i[1819]);
assign l_40[1607]    = ( l_41 [3212] & !i[1819]) | ( l_41 [3213] &  i[1819]);
assign l_40[1608]    = ( l_41 [3214] & !i[1819]) | ( l_41 [3215] &  i[1819]);
assign l_40[1609]    = ( l_41 [3216] & !i[1819]) | ( l_41 [3217] &  i[1819]);
assign l_40[1610]    = ( l_41 [3218] & !i[1819]) | ( l_41 [3219] &  i[1819]);
assign l_40[1611]    = ( l_41 [3220] & !i[1819]) | ( l_41 [3221] &  i[1819]);
assign l_40[1612]    = ( l_41 [3222] & !i[1819]) | ( l_41 [3223] &  i[1819]);
assign l_40[1613]    = ( l_41 [3224] & !i[1819]) | ( l_41 [3225] &  i[1819]);
assign l_40[1614]    = ( l_41 [3226] & !i[1819]) | ( l_41 [3227] &  i[1819]);
assign l_40[1615]    = ( l_41 [3228] & !i[1819]) | ( l_41 [3229] &  i[1819]);
assign l_40[1616]    = ( l_41 [3230] & !i[1819]) | ( l_41 [3231] &  i[1819]);
assign l_40[1617]    = ( l_41 [3232] & !i[1819]) | ( l_41 [3233] &  i[1819]);
assign l_40[1618]    = ( l_41 [3234] & !i[1819]) | ( l_41 [3235] &  i[1819]);
assign l_40[1619]    = ( l_41 [3236] & !i[1819]) | ( l_41 [3237] &  i[1819]);
assign l_40[1620]    = ( l_41 [3238] & !i[1819]) | ( l_41 [3239] &  i[1819]);
assign l_40[1621]    = ( l_41 [3240] & !i[1819]) | ( l_41 [3241] &  i[1819]);
assign l_40[1622]    = ( l_41 [3242] & !i[1819]) | ( l_41 [3243] &  i[1819]);
assign l_40[1623]    = ( l_41 [3244] & !i[1819]) | ( l_41 [3245] &  i[1819]);
assign l_40[1624]    = ( l_41 [3246] & !i[1819]) | ( l_41 [3247] &  i[1819]);
assign l_40[1625]    = ( l_41 [3248] & !i[1819]) | ( l_41 [3249] &  i[1819]);
assign l_40[1626]    = ( l_41 [3250] & !i[1819]) | ( l_41 [3251] &  i[1819]);
assign l_40[1627]    = ( l_41 [3252] & !i[1819]) | ( l_41 [3253] &  i[1819]);
assign l_40[1628]    = ( l_41 [3254] & !i[1819]) | ( l_41 [3255] &  i[1819]);
assign l_40[1629]    = ( l_41 [3256] & !i[1819]) | ( l_41 [3257] &  i[1819]);
assign l_40[1630]    = ( l_41 [3258] & !i[1819]) | ( l_41 [3259] &  i[1819]);
assign l_40[1631]    = ( l_41 [3260] & !i[1819]) | ( l_41 [3261] &  i[1819]);
assign l_40[1632]    = ( l_41 [3262] & !i[1819]) | ( l_41 [3263] &  i[1819]);
assign l_40[1633]    = ( l_41 [3264] & !i[1819]) | ( l_41 [3265] &  i[1819]);
assign l_40[1634]    = ( l_41 [3266] & !i[1819]) | ( l_41 [3267] &  i[1819]);
assign l_40[1635]    = ( l_41 [3268] & !i[1819]) | ( l_41 [3269] &  i[1819]);
assign l_40[1636]    = ( l_41 [3270] & !i[1819]) | ( l_41 [3271] &  i[1819]);
assign l_40[1637]    = ( l_41 [3272] & !i[1819]) | ( l_41 [3273] &  i[1819]);
assign l_40[1638]    = ( l_41 [3274] & !i[1819]) | ( l_41 [3275] &  i[1819]);
assign l_40[1639]    = ( l_41 [3276] & !i[1819]) | ( l_41 [3277] &  i[1819]);
assign l_40[1640]    = ( l_41 [3278] & !i[1819]) | ( l_41 [3279] &  i[1819]);
assign l_40[1641]    = ( l_41 [3280] & !i[1819]) | ( l_41 [3281] &  i[1819]);
assign l_40[1642]    = ( l_41 [3282] & !i[1819]) | ( l_41 [3283] &  i[1819]);
assign l_40[1643]    = ( l_41 [3284] & !i[1819]) | ( l_41 [3285] &  i[1819]);
assign l_40[1644]    = ( l_41 [3286] & !i[1819]) | ( l_41 [3287] &  i[1819]);
assign l_40[1645]    = ( l_41 [3288] & !i[1819]) | ( l_41 [3289] &  i[1819]);
assign l_40[1646]    = ( l_41 [3290] & !i[1819]) | ( l_41 [3291] &  i[1819]);
assign l_40[1647]    = ( l_41 [3292] & !i[1819]) | ( l_41 [3293] &  i[1819]);
assign l_40[1648]    = ( l_41 [3294] & !i[1819]) | ( l_41 [3295] &  i[1819]);
assign l_40[1649]    = ( l_41 [3296] & !i[1819]) | ( l_41 [3297] &  i[1819]);
assign l_40[1650]    = ( l_41 [3298] & !i[1819]) | ( l_41 [3299] &  i[1819]);
assign l_40[1651]    = ( l_41 [3300] & !i[1819]) | ( l_41 [3301] &  i[1819]);
assign l_40[1652]    = ( l_41 [3302] & !i[1819]) | ( l_41 [3303] &  i[1819]);
assign l_40[1653]    = ( l_41 [3304] & !i[1819]) | ( l_41 [3305] &  i[1819]);
assign l_40[1654]    = ( l_41 [3306] & !i[1819]) | ( l_41 [3307] &  i[1819]);
assign l_40[1655]    = ( l_41 [3308] & !i[1819]) | ( l_41 [3309] &  i[1819]);
assign l_40[1656]    = ( l_41 [3310] & !i[1819]) | ( l_41 [3311] &  i[1819]);
assign l_40[1657]    = ( l_41 [3312] & !i[1819]) | ( l_41 [3313] &  i[1819]);
assign l_40[1658]    = ( l_41 [3314] & !i[1819]) | ( l_41 [3315] &  i[1819]);
assign l_40[1659]    = ( l_41 [3316] & !i[1819]) | ( l_41 [3317] &  i[1819]);
assign l_40[1660]    = ( l_41 [3318] & !i[1819]) | ( l_41 [3319] &  i[1819]);
assign l_40[1661]    = ( l_41 [3320] & !i[1819]) | ( l_41 [3321] &  i[1819]);
assign l_40[1662]    = ( l_41 [3322] & !i[1819]) | ( l_41 [3323] &  i[1819]);
assign l_40[1663]    = ( l_41 [3324] & !i[1819]) | ( l_41 [3325] &  i[1819]);
assign l_40[1664]    = ( l_41 [3326] & !i[1819]) | ( l_41 [3327] &  i[1819]);
assign l_40[1665]    = ( l_41 [3328] & !i[1819]) | ( l_41 [3329] &  i[1819]);
assign l_40[1666]    = ( l_41 [3330] & !i[1819]) | ( l_41 [3331] &  i[1819]);
assign l_40[1667]    = ( l_41 [3332] & !i[1819]) | ( l_41 [3333] &  i[1819]);
assign l_40[1668]    = ( l_41 [3334] & !i[1819]) | ( l_41 [3335] &  i[1819]);
assign l_40[1669]    = ( l_41 [3336] & !i[1819]) | ( l_41 [3337] &  i[1819]);
assign l_40[1670]    = ( l_41 [3338] & !i[1819]) | ( l_41 [3339] &  i[1819]);
assign l_40[1671]    = ( l_41 [3340] & !i[1819]) | ( l_41 [3341] &  i[1819]);
assign l_40[1672]    = ( l_41 [3342] & !i[1819]) | ( l_41 [3343] &  i[1819]);
assign l_40[1673]    = ( l_41 [3344] & !i[1819]) | ( l_41 [3345] &  i[1819]);
assign l_40[1674]    = ( l_41 [3346] & !i[1819]) | ( l_41 [3347] &  i[1819]);
assign l_40[1675]    = ( l_41 [3348] & !i[1819]) | ( l_41 [3349] &  i[1819]);
assign l_40[1676]    = ( l_41 [3350] & !i[1819]) | ( l_41 [3351] &  i[1819]);
assign l_40[1677]    = ( l_41 [3352] & !i[1819]) | ( l_41 [3353] &  i[1819]);
assign l_40[1678]    = ( l_41 [3354] & !i[1819]) | ( l_41 [3355] &  i[1819]);
assign l_40[1679]    = ( l_41 [3356] & !i[1819]) | ( l_41 [3357] &  i[1819]);
assign l_40[1680]    = ( l_41 [3358] & !i[1819]) | ( l_41 [3359] &  i[1819]);
assign l_40[1681]    = ( l_41 [3360] & !i[1819]) | ( l_41 [3361] &  i[1819]);
assign l_40[1682]    = ( l_41 [3362] & !i[1819]) | ( l_41 [3363] &  i[1819]);
assign l_40[1683]    = ( l_41 [3364] & !i[1819]) | ( l_41 [3365] &  i[1819]);
assign l_40[1684]    = ( l_41 [3366] & !i[1819]) | ( l_41 [3367] &  i[1819]);
assign l_40[1685]    = ( l_41 [3368] & !i[1819]) | ( l_41 [3369] &  i[1819]);
assign l_40[1686]    = ( l_41 [3370] & !i[1819]) | ( l_41 [3371] &  i[1819]);
assign l_40[1687]    = ( l_41 [3372] & !i[1819]) | ( l_41 [3373] &  i[1819]);
assign l_40[1688]    = ( l_41 [3374] & !i[1819]) | ( l_41 [3375] &  i[1819]);
assign l_40[1689]    = ( l_41 [3376] & !i[1819]) | ( l_41 [3377] &  i[1819]);
assign l_40[1690]    = ( l_41 [3378] & !i[1819]) | ( l_41 [3379] &  i[1819]);
assign l_40[1691]    = ( l_41 [3380] & !i[1819]) | ( l_41 [3381] &  i[1819]);
assign l_40[1692]    = ( l_41 [3382] & !i[1819]) | ( l_41 [3383] &  i[1819]);
assign l_40[1693]    = ( l_41 [3384] & !i[1819]) | ( l_41 [3385] &  i[1819]);
assign l_40[1694]    = ( l_41 [3386] & !i[1819]) | ( l_41 [3387] &  i[1819]);
assign l_40[1695]    = ( l_41 [3388] & !i[1819]) | ( l_41 [3389] &  i[1819]);
assign l_40[1696]    = ( l_41 [3390] & !i[1819]) | ( l_41 [3391] &  i[1819]);
assign l_40[1697]    = ( l_41 [3392] & !i[1819]) | ( l_41 [3393] &  i[1819]);
assign l_40[1698]    = ( l_41 [3394] & !i[1819]) | ( l_41 [3395] &  i[1819]);
assign l_40[1699]    = ( l_41 [3396] & !i[1819]) | ( l_41 [3397] &  i[1819]);
assign l_40[1700]    = ( l_41 [3398] & !i[1819]) | ( l_41 [3399] &  i[1819]);
assign l_40[1701]    = ( l_41 [3400] & !i[1819]) | ( l_41 [3401] &  i[1819]);
assign l_40[1702]    = ( l_41 [3402] & !i[1819]) | ( l_41 [3403] &  i[1819]);
assign l_40[1703]    = ( l_41 [3404] & !i[1819]) | ( l_41 [3405] &  i[1819]);
assign l_40[1704]    = ( l_41 [3406] & !i[1819]) | ( l_41 [3407] &  i[1819]);
assign l_40[1705]    = ( l_41 [3408] & !i[1819]) | ( l_41 [3409] &  i[1819]);
assign l_40[1706]    = ( l_41 [3410] & !i[1819]) | ( l_41 [3411] &  i[1819]);
assign l_40[1707]    = ( l_41 [3412] & !i[1819]) | ( l_41 [3413] &  i[1819]);
assign l_40[1708]    = ( l_41 [3414] & !i[1819]) | ( l_41 [3415] &  i[1819]);
assign l_40[1709]    = ( l_41 [3416] & !i[1819]) | ( l_41 [3417] &  i[1819]);
assign l_40[1710]    = ( l_41 [3418] & !i[1819]) | ( l_41 [3419] &  i[1819]);
assign l_40[1711]    = ( l_41 [3420] & !i[1819]) | ( l_41 [3421] &  i[1819]);
assign l_40[1712]    = ( l_41 [3422] & !i[1819]) | ( l_41 [3423] &  i[1819]);
assign l_40[1713]    = ( l_41 [3424] & !i[1819]) | ( l_41 [3425] &  i[1819]);
assign l_40[1714]    = ( l_41 [3426] & !i[1819]) | ( l_41 [3427] &  i[1819]);
assign l_40[1715]    = ( l_41 [3428] & !i[1819]) | ( l_41 [3429] &  i[1819]);
assign l_40[1716]    = ( l_41 [3430] & !i[1819]) | ( l_41 [3431] &  i[1819]);
assign l_40[1717]    = ( l_41 [3432] & !i[1819]) | ( l_41 [3433] &  i[1819]);
assign l_40[1718]    = ( l_41 [3434] & !i[1819]) | ( l_41 [3435] &  i[1819]);
assign l_40[1719]    = ( l_41 [3436] & !i[1819]) | ( l_41 [3437] &  i[1819]);
assign l_40[1720]    = ( l_41 [3438] & !i[1819]) | ( l_41 [3439] &  i[1819]);
assign l_40[1721]    = ( l_41 [3440] & !i[1819]) | ( l_41 [3441] &  i[1819]);
assign l_40[1722]    = ( l_41 [3442] & !i[1819]) | ( l_41 [3443] &  i[1819]);
assign l_40[1723]    = ( l_41 [3444] & !i[1819]) | ( l_41 [3445] &  i[1819]);
assign l_40[1724]    = ( l_41 [3446] & !i[1819]) | ( l_41 [3447] &  i[1819]);
assign l_40[1725]    = ( l_41 [3448] & !i[1819]) | ( l_41 [3449] &  i[1819]);
assign l_40[1726]    = ( l_41 [3450] & !i[1819]) | ( l_41 [3451] &  i[1819]);
assign l_40[1727]    = ( l_41 [3452] & !i[1819]) | ( l_41 [3453] &  i[1819]);
assign l_40[1728]    = ( l_41 [3454] & !i[1819]) | ( l_41 [3455] &  i[1819]);
assign l_40[1729]    = ( l_41 [3456] & !i[1819]) | ( l_41 [3457] &  i[1819]);
assign l_40[1730]    = ( l_41 [3458] & !i[1819]) | ( l_41 [3459] &  i[1819]);
assign l_40[1731]    = ( l_41 [3460] & !i[1819]) | ( l_41 [3461] &  i[1819]);
assign l_40[1732]    = ( l_41 [3462] & !i[1819]) | ( l_41 [3463] &  i[1819]);
assign l_40[1733]    = ( l_41 [3464] & !i[1819]) | ( l_41 [3465] &  i[1819]);
assign l_40[1734]    = ( l_41 [3466] & !i[1819]) | ( l_41 [3467] &  i[1819]);
assign l_40[1735]    = ( l_41 [3468] & !i[1819]) | ( l_41 [3469] &  i[1819]);
assign l_40[1736]    = ( l_41 [3470] & !i[1819]) | ( l_41 [3471] &  i[1819]);
assign l_40[1737]    = ( l_41 [3472] & !i[1819]) | ( l_41 [3473] &  i[1819]);
assign l_40[1738]    = ( l_41 [3474] & !i[1819]) | ( l_41 [3475] &  i[1819]);
assign l_40[1739]    = ( l_41 [3476] & !i[1819]) | ( l_41 [3477] &  i[1819]);
assign l_40[1740]    = ( l_41 [3478] & !i[1819]) | ( l_41 [3479] &  i[1819]);
assign l_40[1741]    = ( l_41 [3480] & !i[1819]) | ( l_41 [3481] &  i[1819]);
assign l_40[1742]    = ( l_41 [3482] & !i[1819]) | ( l_41 [3483] &  i[1819]);
assign l_40[1743]    = ( l_41 [3484] & !i[1819]) | ( l_41 [3485] &  i[1819]);
assign l_40[1744]    = ( l_41 [3486] & !i[1819]) | ( l_41 [3487] &  i[1819]);
assign l_40[1745]    = ( l_41 [3488] & !i[1819]) | ( l_41 [3489] &  i[1819]);
assign l_40[1746]    = ( l_41 [3490] & !i[1819]) | ( l_41 [3491] &  i[1819]);
assign l_40[1747]    = ( l_41 [3492] & !i[1819]) | ( l_41 [3493] &  i[1819]);
assign l_40[1748]    = ( l_41 [3494] & !i[1819]) | ( l_41 [3495] &  i[1819]);
assign l_40[1749]    = ( l_41 [3496] & !i[1819]) | ( l_41 [3497] &  i[1819]);
assign l_40[1750]    = ( l_41 [3498] & !i[1819]) | ( l_41 [3499] &  i[1819]);
assign l_40[1751]    = ( l_41 [3500] & !i[1819]) | ( l_41 [3501] &  i[1819]);
assign l_40[1752]    = ( l_41 [3502] & !i[1819]) | ( l_41 [3503] &  i[1819]);
assign l_40[1753]    = ( l_41 [3504] & !i[1819]) | ( l_41 [3505] &  i[1819]);
assign l_40[1754]    = ( l_41 [3506] & !i[1819]) | ( l_41 [3507] &  i[1819]);
assign l_40[1755]    = ( l_41 [3508] & !i[1819]) | ( l_41 [3509] &  i[1819]);
assign l_40[1756]    = ( l_41 [3510] & !i[1819]) | ( l_41 [3511] &  i[1819]);
assign l_40[1757]    = ( l_41 [3512] & !i[1819]) | ( l_41 [3513] &  i[1819]);
assign l_40[1758]    = ( l_41 [3514] & !i[1819]) | ( l_41 [3515] &  i[1819]);
assign l_40[1759]    = ( l_41 [3516] & !i[1819]) | ( l_41 [3517] &  i[1819]);
assign l_40[1760]    = ( l_41 [3518] & !i[1819]) | ( l_41 [3519] &  i[1819]);
assign l_40[1761]    = ( l_41 [3520] & !i[1819]) | ( l_41 [3521] &  i[1819]);
assign l_40[1762]    = ( l_41 [3522] & !i[1819]) | ( l_41 [3523] &  i[1819]);
assign l_40[1763]    = ( l_41 [3524] & !i[1819]) | ( l_41 [3525] &  i[1819]);
assign l_40[1764]    = ( l_41 [3526] & !i[1819]) | ( l_41 [3527] &  i[1819]);
assign l_40[1765]    = ( l_41 [3528] & !i[1819]) | ( l_41 [3529] &  i[1819]);
assign l_40[1766]    = ( l_41 [3530] & !i[1819]) | ( l_41 [3531] &  i[1819]);
assign l_40[1767]    = ( l_41 [3532] & !i[1819]) | ( l_41 [3533] &  i[1819]);
assign l_40[1768]    = ( l_41 [3534] & !i[1819]) | ( l_41 [3535] &  i[1819]);
assign l_40[1769]    = ( l_41 [3536] & !i[1819]) | ( l_41 [3537] &  i[1819]);
assign l_40[1770]    = ( l_41 [3538] & !i[1819]) | ( l_41 [3539] &  i[1819]);
assign l_40[1771]    = ( l_41 [3540] & !i[1819]) | ( l_41 [3541] &  i[1819]);
assign l_40[1772]    = ( l_41 [3542] & !i[1819]) | ( l_41 [3543] &  i[1819]);
assign l_40[1773]    = ( l_41 [3544] & !i[1819]) | ( l_41 [3545] &  i[1819]);
assign l_40[1774]    = ( l_41 [3546] & !i[1819]) | ( l_41 [3547] &  i[1819]);
assign l_40[1775]    = ( l_41 [3548] & !i[1819]) | ( l_41 [3549] &  i[1819]);
assign l_40[1776]    = ( l_41 [3550] & !i[1819]) | ( l_41 [3551] &  i[1819]);
assign l_40[1777]    = ( l_41 [3552] & !i[1819]) | ( l_41 [3553] &  i[1819]);
assign l_40[1778]    = ( l_41 [3554] & !i[1819]) | ( l_41 [3555] &  i[1819]);
assign l_40[1779]    = ( l_41 [3556] & !i[1819]) | ( l_41 [3557] &  i[1819]);
assign l_40[1780]    = ( l_41 [3558] & !i[1819]) | ( l_41 [3559] &  i[1819]);
assign l_40[1781]    = ( l_41 [3560] & !i[1819]) | ( l_41 [3561] &  i[1819]);
assign l_40[1782]    = ( l_41 [3562] & !i[1819]) | ( l_41 [3563] &  i[1819]);
assign l_40[1783]    = ( l_41 [3564] & !i[1819]) | ( l_41 [3565] &  i[1819]);
assign l_40[1784]    = ( l_41 [3566] & !i[1819]) | ( l_41 [3567] &  i[1819]);
assign l_40[1785]    = ( l_41 [3568] & !i[1819]) | ( l_41 [3569] &  i[1819]);
assign l_40[1786]    = ( l_41 [3570] & !i[1819]) | ( l_41 [3571] &  i[1819]);
assign l_40[1787]    = ( l_41 [3572] & !i[1819]) | ( l_41 [3573] &  i[1819]);
assign l_40[1788]    = ( l_41 [3574] & !i[1819]) | ( l_41 [3575] &  i[1819]);
assign l_40[1789]    = ( l_41 [3576] & !i[1819]) | ( l_41 [3577] &  i[1819]);
assign l_40[1790]    = ( l_41 [3578] & !i[1819]) | ( l_41 [3579] &  i[1819]);
assign l_40[1791]    = ( l_41 [3580] & !i[1819]) | ( l_41 [3581] &  i[1819]);
assign l_40[1792]    = ( l_41 [3582] & !i[1819]) | ( l_41 [3583] &  i[1819]);
assign l_40[1793]    = ( l_41 [3584] & !i[1819]) | ( l_41 [3585] &  i[1819]);
assign l_40[1794]    = ( l_41 [3586] & !i[1819]) | ( l_41 [3587] &  i[1819]);
assign l_40[1795]    = ( l_41 [3588] & !i[1819]) | ( l_41 [3589] &  i[1819]);
assign l_40[1796]    = ( l_41 [3590] & !i[1819]) | ( l_41 [3591] &  i[1819]);
assign l_40[1797]    = ( l_41 [3592] & !i[1819]) | ( l_41 [3593] &  i[1819]);
assign l_40[1798]    = ( l_41 [3594] & !i[1819]) | ( l_41 [3595] &  i[1819]);
assign l_40[1799]    = ( l_41 [3596] & !i[1819]) | ( l_41 [3597] &  i[1819]);
assign l_40[1800]    = ( l_41 [3598] & !i[1819]) | ( l_41 [3599] &  i[1819]);
assign l_40[1801]    = ( l_41 [3600] & !i[1819]) | ( l_41 [3601] &  i[1819]);
assign l_40[1802]    = ( l_41 [3602] & !i[1819]) | ( l_41 [3603] &  i[1819]);
assign l_40[1803]    = ( l_41 [3604] & !i[1819]) | ( l_41 [3605] &  i[1819]);
assign l_40[1804]    = ( l_41 [3606] & !i[1819]) | ( l_41 [3607] &  i[1819]);
assign l_40[1805]    = ( l_41 [3608] & !i[1819]) | ( l_41 [3609] &  i[1819]);
assign l_40[1806]    = ( l_41 [3610] & !i[1819]) | ( l_41 [3611] &  i[1819]);
assign l_40[1807]    = ( l_41 [3612] & !i[1819]) | ( l_41 [3613] &  i[1819]);
assign l_40[1808]    = ( l_41 [3614] & !i[1819]) | ( l_41 [3615] &  i[1819]);
assign l_40[1809]    = ( l_41 [3616] & !i[1819]) | ( l_41 [3617] &  i[1819]);
assign l_40[1810]    = ( l_41 [3618] & !i[1819]) | ( l_41 [3619] &  i[1819]);
assign l_40[1811]    = ( l_41 [3620] & !i[1819]) | ( l_41 [3621] &  i[1819]);
assign l_40[1812]    = ( l_41 [3622] & !i[1819]) | ( l_41 [3623] &  i[1819]);
assign l_40[1813]    = ( l_41 [3624] & !i[1819]) | ( l_41 [3625] &  i[1819]);
assign l_40[1814]    = ( l_41 [3626] & !i[1819]) | ( l_41 [3627] &  i[1819]);
assign l_40[1815]    = ( l_41 [3628] & !i[1819]) | ( l_41 [3629] &  i[1819]);
assign l_40[1816]    = ( l_41 [3630] & !i[1819]) | ( l_41 [3631] &  i[1819]);
assign l_40[1817]    = ( l_41 [3632] & !i[1819]) | ( l_41 [3633] &  i[1819]);
assign l_40[1818]    = ( l_41 [3634] & !i[1819]) | ( l_41 [3635] &  i[1819]);
assign l_40[1819]    = ( l_41 [3636] & !i[1819]) | ( l_41 [3637] &  i[1819]);
assign l_40[1820]    = ( l_41 [3638] & !i[1819]) | ( l_41 [3639] &  i[1819]);
assign l_40[1821]    = ( l_41 [3640] & !i[1819]) | ( l_41 [3641] &  i[1819]);
assign l_40[1822]    = ( l_41 [3642] & !i[1819]) | ( l_41 [3643] &  i[1819]);
assign l_40[1823]    = ( l_41 [3644] & !i[1819]) | ( l_41 [3645] &  i[1819]);
assign l_40[1824]    = ( l_41 [3646] & !i[1819]) | ( l_41 [3647] &  i[1819]);
assign l_40[1825]    = ( l_41 [3648] & !i[1819]) | ( l_41 [3649] &  i[1819]);
assign l_40[1826]    = ( l_41 [3650] & !i[1819]) | ( l_41 [3651] &  i[1819]);
assign l_40[1827]    = ( l_41 [3652] & !i[1819]) | ( l_41 [3653] &  i[1819]);
assign l_40[1828]    = ( l_41 [3654] & !i[1819]) | ( l_41 [3655] &  i[1819]);
assign l_40[1829]    = ( l_41 [3656] & !i[1819]) | ( l_41 [3657] &  i[1819]);
assign l_40[1830]    = ( l_41 [3658] & !i[1819]) | ( l_41 [3659] &  i[1819]);
assign l_40[1831]    = ( l_41 [3660] & !i[1819]) | ( l_41 [3661] &  i[1819]);
assign l_40[1832]    = ( l_41 [3662] & !i[1819]) | ( l_41 [3663] &  i[1819]);
assign l_40[1833]    = ( l_41 [3664] & !i[1819]) | ( l_41 [3665] &  i[1819]);
assign l_40[1834]    = ( l_41 [3666] & !i[1819]) | ( l_41 [3667] &  i[1819]);
assign l_40[1835]    = ( l_41 [3668] & !i[1819]) | ( l_41 [3669] &  i[1819]);
assign l_40[1836]    = ( l_41 [3670] & !i[1819]) | ( l_41 [3671] &  i[1819]);
assign l_40[1837]    = ( l_41 [3672] & !i[1819]) | ( l_41 [3673] &  i[1819]);
assign l_40[1838]    = ( l_41 [3674] & !i[1819]) | ( l_41 [3675] &  i[1819]);
assign l_40[1839]    = ( l_41 [3676] & !i[1819]) | ( l_41 [3677] &  i[1819]);
assign l_40[1840]    = ( l_41 [3678] & !i[1819]) | ( l_41 [3679] &  i[1819]);
assign l_40[1841]    = ( l_41 [3680] & !i[1819]) | ( l_41 [3681] &  i[1819]);
assign l_40[1842]    = ( l_41 [3682] & !i[1819]) | ( l_41 [3683] &  i[1819]);
assign l_40[1843]    = ( l_41 [3684] & !i[1819]) | ( l_41 [3685] &  i[1819]);
assign l_40[1844]    = ( l_41 [3686] & !i[1819]) | ( l_41 [3687] &  i[1819]);
assign l_40[1845]    = ( l_41 [3688] & !i[1819]) | ( l_41 [3689] &  i[1819]);
assign l_40[1846]    = ( l_41 [3690] & !i[1819]) | ( l_41 [3691] &  i[1819]);
assign l_40[1847]    = ( l_41 [3692] & !i[1819]) | ( l_41 [3693] &  i[1819]);
assign l_40[1848]    = ( l_41 [3694] & !i[1819]) | ( l_41 [3695] &  i[1819]);
assign l_40[1849]    = ( l_41 [3696] & !i[1819]) | ( l_41 [3697] &  i[1819]);
assign l_40[1850]    = ( l_41 [3698] & !i[1819]) | ( l_41 [3699] &  i[1819]);
assign l_40[1851]    = ( l_41 [3700] & !i[1819]) | ( l_41 [3701] &  i[1819]);
assign l_40[1852]    = ( l_41 [3702] & !i[1819]) | ( l_41 [3703] &  i[1819]);
assign l_40[1853]    = ( l_41 [3704] & !i[1819]) | ( l_41 [3705] &  i[1819]);
assign l_40[1854]    = ( l_41 [3706] & !i[1819]) | ( l_41 [3707] &  i[1819]);
assign l_40[1855]    = ( l_41 [3708] & !i[1819]) | ( l_41 [3709] &  i[1819]);
assign l_40[1856]    = ( l_41 [3710] & !i[1819]) | ( l_41 [3711] &  i[1819]);
assign l_40[1857]    = ( l_41 [3712] & !i[1819]) | ( l_41 [3713] &  i[1819]);
assign l_40[1858]    = ( l_41 [3714] & !i[1819]) | ( l_41 [3715] &  i[1819]);
assign l_40[1859]    = ( l_41 [3716] & !i[1819]) | ( l_41 [3717] &  i[1819]);
assign l_40[1860]    = ( l_41 [3718] & !i[1819]) | ( l_41 [3719] &  i[1819]);
assign l_40[1861]    = ( l_41 [3720] & !i[1819]) | ( l_41 [3721] &  i[1819]);
assign l_40[1862]    = ( l_41 [3722] & !i[1819]) | ( l_41 [3723] &  i[1819]);
assign l_40[1863]    = ( l_41 [3724] & !i[1819]) | ( l_41 [3725] &  i[1819]);
assign l_40[1864]    = ( l_41 [3726] & !i[1819]) | ( l_41 [3727] &  i[1819]);
assign l_40[1865]    = ( l_41 [3728] & !i[1819]) | ( l_41 [3729] &  i[1819]);
assign l_40[1866]    = ( l_41 [3730] & !i[1819]) | ( l_41 [3731] &  i[1819]);
assign l_40[1867]    = ( l_41 [3732] & !i[1819]) | ( l_41 [3733] &  i[1819]);
assign l_40[1868]    = ( l_41 [3734] & !i[1819]) | ( l_41 [3735] &  i[1819]);
assign l_40[1869]    = ( l_41 [3736] & !i[1819]) | ( l_41 [3737] &  i[1819]);
assign l_40[1870]    = ( l_41 [3738] & !i[1819]) | ( l_41 [3739] &  i[1819]);
assign l_40[1871]    = ( l_41 [3740] & !i[1819]) | ( l_41 [3741] &  i[1819]);
assign l_40[1872]    = ( l_41 [3742] & !i[1819]) | ( l_41 [3743] &  i[1819]);
assign l_40[1873]    = ( l_41 [3744] & !i[1819]) | ( l_41 [3745] &  i[1819]);
assign l_40[1874]    = ( l_41 [3746] & !i[1819]) | ( l_41 [3747] &  i[1819]);
assign l_40[1875]    = ( l_41 [3748] & !i[1819]) | ( l_41 [3749] &  i[1819]);
assign l_40[1876]    = ( l_41 [3750] & !i[1819]) | ( l_41 [3751] &  i[1819]);
assign l_40[1877]    = ( l_41 [3752] & !i[1819]) | ( l_41 [3753] &  i[1819]);
assign l_40[1878]    = ( l_41 [3754] & !i[1819]) | ( l_41 [3755] &  i[1819]);
assign l_40[1879]    = ( l_41 [3756] & !i[1819]) | ( l_41 [3757] &  i[1819]);
assign l_40[1880]    = ( l_41 [3758] & !i[1819]) | ( l_41 [3759] &  i[1819]);
assign l_40[1881]    = ( l_41 [3760] & !i[1819]) | ( l_41 [3761] &  i[1819]);
assign l_40[1882]    = ( l_41 [3762] & !i[1819]) | ( l_41 [3763] &  i[1819]);
assign l_40[1883]    = ( l_41 [3764] & !i[1819]) | ( l_41 [3765] &  i[1819]);
assign l_40[1884]    = ( l_41 [3766] & !i[1819]) | ( l_41 [3767] &  i[1819]);
assign l_40[1885]    = ( l_41 [3768] & !i[1819]) | ( l_41 [3769] &  i[1819]);
assign l_40[1886]    = ( l_41 [3770] & !i[1819]) | ( l_41 [3771] &  i[1819]);
assign l_40[1887]    = ( l_41 [3772] & !i[1819]) | ( l_41 [3773] &  i[1819]);
assign l_40[1888]    = ( l_41 [3774] & !i[1819]) | ( l_41 [3775] &  i[1819]);
assign l_40[1889]    = ( l_41 [3776] & !i[1819]) | ( l_41 [3777] &  i[1819]);
assign l_40[1890]    = ( l_41 [3778] & !i[1819]) | ( l_41 [3779] &  i[1819]);
assign l_40[1891]    = ( l_41 [3780] & !i[1819]) | ( l_41 [3781] &  i[1819]);
assign l_40[1892]    = ( l_41 [3782] & !i[1819]) | ( l_41 [3783] &  i[1819]);
assign l_40[1893]    = ( l_41 [3784] & !i[1819]) | ( l_41 [3785] &  i[1819]);
assign l_40[1894]    = ( l_41 [3786] & !i[1819]) | ( l_41 [3787] &  i[1819]);
assign l_40[1895]    = ( l_41 [3788] & !i[1819]) | ( l_41 [3789] &  i[1819]);
assign l_40[1896]    = ( l_41 [3790] & !i[1819]) | ( l_41 [3791] &  i[1819]);
assign l_40[1897]    = ( l_41 [3792] & !i[1819]) | ( l_41 [3793] &  i[1819]);
assign l_40[1898]    = ( l_41 [3794] & !i[1819]) | ( l_41 [3795] &  i[1819]);
assign l_40[1899]    = ( l_41 [3796] & !i[1819]) | ( l_41 [3797] &  i[1819]);
assign l_40[1900]    = ( l_41 [3798] & !i[1819]) | ( l_41 [3799] &  i[1819]);
assign l_40[1901]    = ( l_41 [3800] & !i[1819]) | ( l_41 [3801] &  i[1819]);
assign l_40[1902]    = ( l_41 [3802] & !i[1819]) | ( l_41 [3803] &  i[1819]);
assign l_40[1903]    = ( l_41 [3804] & !i[1819]) | ( l_41 [3805] &  i[1819]);
assign l_40[1904]    = ( l_41 [3806] & !i[1819]) | ( l_41 [3807] &  i[1819]);
assign l_40[1905]    = ( l_41 [3808] & !i[1819]) | ( l_41 [3809] &  i[1819]);
assign l_40[1906]    = ( l_41 [3810] & !i[1819]) | ( l_41 [3811] &  i[1819]);
assign l_40[1907]    = ( l_41 [3812] & !i[1819]) | ( l_41 [3813] &  i[1819]);
assign l_40[1908]    = ( l_41 [3814] & !i[1819]) | ( l_41 [3815] &  i[1819]);
assign l_40[1909]    = ( l_41 [3816] & !i[1819]) | ( l_41 [3817] &  i[1819]);
assign l_40[1910]    = ( l_41 [3818] & !i[1819]) | ( l_41 [3819] &  i[1819]);
assign l_40[1911]    = ( l_41 [3820] & !i[1819]) | ( l_41 [3821] &  i[1819]);
assign l_40[1912]    = ( l_41 [3822] & !i[1819]) | ( l_41 [3823] &  i[1819]);
assign l_40[1913]    = ( l_41 [3824] & !i[1819]) | ( l_41 [3825] &  i[1819]);
assign l_40[1914]    = ( l_41 [3826] & !i[1819]) | ( l_41 [3827] &  i[1819]);
assign l_40[1915]    = ( l_41 [3828] & !i[1819]) | ( l_41 [3829] &  i[1819]);
assign l_40[1916]    = ( l_41 [3830] & !i[1819]) | ( l_41 [3831] &  i[1819]);
assign l_40[1917]    = ( l_41 [3832] & !i[1819]) | ( l_41 [3833] &  i[1819]);
assign l_40[1918]    = ( l_41 [3834] & !i[1819]) | ( l_41 [3835] &  i[1819]);
assign l_40[1919]    = ( l_41 [3836] & !i[1819]) | ( l_41 [3837] &  i[1819]);
assign l_40[1920]    = ( l_41 [3838] & !i[1819]) | ( l_41 [3839] &  i[1819]);
assign l_40[1921]    = ( l_41 [3840] & !i[1819]) | ( l_41 [3841] &  i[1819]);
assign l_40[1922]    = ( l_41 [3842] & !i[1819]) | ( l_41 [3843] &  i[1819]);
assign l_40[1923]    = ( l_41 [3844] & !i[1819]) | ( l_41 [3845] &  i[1819]);
assign l_40[1924]    = ( l_41 [3846] & !i[1819]) | ( l_41 [3847] &  i[1819]);
assign l_40[1925]    = ( l_41 [3848] & !i[1819]) | ( l_41 [3849] &  i[1819]);
assign l_40[1926]    = ( l_41 [3850] & !i[1819]) | ( l_41 [3851] &  i[1819]);
assign l_40[1927]    = ( l_41 [3852] & !i[1819]) | ( l_41 [3853] &  i[1819]);
assign l_40[1928]    = ( l_41 [3854] & !i[1819]) | ( l_41 [3855] &  i[1819]);
assign l_40[1929]    = ( l_41 [3856] & !i[1819]) | ( l_41 [3857] &  i[1819]);
assign l_40[1930]    = ( l_41 [3858] & !i[1819]) | ( l_41 [3859] &  i[1819]);
assign l_40[1931]    = ( l_41 [3860] & !i[1819]) | ( l_41 [3861] &  i[1819]);
assign l_40[1932]    = ( l_41 [3862] & !i[1819]) | ( l_41 [3863] &  i[1819]);
assign l_40[1933]    = ( l_41 [3864] & !i[1819]) | ( l_41 [3865] &  i[1819]);
assign l_40[1934]    = ( l_41 [3866] & !i[1819]) | ( l_41 [3867] &  i[1819]);
assign l_40[1935]    = ( l_41 [3868] & !i[1819]) | ( l_41 [3869] &  i[1819]);
assign l_40[1936]    = ( l_41 [3870] & !i[1819]) | ( l_41 [3871] &  i[1819]);
assign l_40[1937]    = ( l_41 [3872] & !i[1819]) | ( l_41 [3873] &  i[1819]);
assign l_40[1938]    = ( l_41 [3874] & !i[1819]) | ( l_41 [3875] &  i[1819]);
assign l_40[1939]    = ( l_41 [3876] & !i[1819]) | ( l_41 [3877] &  i[1819]);
assign l_40[1940]    = ( l_41 [3878] & !i[1819]) | ( l_41 [3879] &  i[1819]);
assign l_40[1941]    = ( l_41 [3880] & !i[1819]) | ( l_41 [3881] &  i[1819]);
assign l_40[1942]    = ( l_41 [3882] & !i[1819]) | ( l_41 [3883] &  i[1819]);
assign l_40[1943]    = ( l_41 [3884] & !i[1819]) | ( l_41 [3885] &  i[1819]);
assign l_40[1944]    = ( l_41 [3886] & !i[1819]) | ( l_41 [3887] &  i[1819]);
assign l_40[1945]    = ( l_41 [3888] & !i[1819]) | ( l_41 [3889] &  i[1819]);
assign l_40[1946]    = ( l_41 [3890] & !i[1819]) | ( l_41 [3891] &  i[1819]);
assign l_40[1947]    = ( l_41 [3892] & !i[1819]) | ( l_41 [3893] &  i[1819]);
assign l_40[1948]    = ( l_41 [3894] & !i[1819]) | ( l_41 [3895] &  i[1819]);
assign l_40[1949]    = ( l_41 [3896] & !i[1819]) | ( l_41 [3897] &  i[1819]);
assign l_40[1950]    = ( l_41 [3898] & !i[1819]) | ( l_41 [3899] &  i[1819]);
assign l_40[1951]    = ( l_41 [3900] & !i[1819]) | ( l_41 [3901] &  i[1819]);
assign l_40[1952]    = ( l_41 [3902] & !i[1819]) | ( l_41 [3903] &  i[1819]);
assign l_40[1953]    = ( l_41 [3904] & !i[1819]) | ( l_41 [3905] &  i[1819]);
assign l_40[1954]    = ( l_41 [3906] & !i[1819]) | ( l_41 [3907] &  i[1819]);
assign l_40[1955]    = ( l_41 [3908] & !i[1819]) | ( l_41 [3909] &  i[1819]);
assign l_40[1956]    = ( l_41 [3910] & !i[1819]) | ( l_41 [3911] &  i[1819]);
assign l_40[1957]    = ( l_41 [3912] & !i[1819]) | ( l_41 [3913] &  i[1819]);
assign l_40[1958]    = ( l_41 [3914] & !i[1819]) | ( l_41 [3915] &  i[1819]);
assign l_40[1959]    = ( l_41 [3916] & !i[1819]) | ( l_41 [3917] &  i[1819]);
assign l_40[1960]    = ( l_41 [3918] & !i[1819]) | ( l_41 [3919] &  i[1819]);
assign l_40[1961]    = ( l_41 [3920] & !i[1819]) | ( l_41 [3921] &  i[1819]);
assign l_40[1962]    = ( l_41 [3922] & !i[1819]) | ( l_41 [3923] &  i[1819]);
assign l_40[1963]    = ( l_41 [3924] & !i[1819]) | ( l_41 [3925] &  i[1819]);
assign l_40[1964]    = ( l_41 [3926] & !i[1819]) | ( l_41 [3927] &  i[1819]);
assign l_40[1965]    = ( l_41 [3928] & !i[1819]) | ( l_41 [3929] &  i[1819]);
assign l_40[1966]    = ( l_41 [3930] & !i[1819]) | ( l_41 [3931] &  i[1819]);
assign l_40[1967]    = ( l_41 [3932] & !i[1819]) | ( l_41 [3933] &  i[1819]);
assign l_40[1968]    = ( l_41 [3934] & !i[1819]) | ( l_41 [3935] &  i[1819]);
assign l_40[1969]    = ( l_41 [3936] & !i[1819]) | ( l_41 [3937] &  i[1819]);
assign l_40[1970]    = ( l_41 [3938] & !i[1819]) | ( l_41 [3939] &  i[1819]);
assign l_40[1971]    = ( l_41 [3940] & !i[1819]) | ( l_41 [3941] &  i[1819]);
assign l_40[1972]    = ( l_41 [3942] & !i[1819]) | ( l_41 [3943] &  i[1819]);
assign l_40[1973]    = ( l_41 [3944] & !i[1819]) | ( l_41 [3945] &  i[1819]);
assign l_40[1974]    = ( l_41 [3946] & !i[1819]) | ( l_41 [3947] &  i[1819]);
assign l_40[1975]    = ( l_41 [3948] & !i[1819]) | ( l_41 [3949] &  i[1819]);
assign l_40[1976]    = ( l_41 [3950] & !i[1819]) | ( l_41 [3951] &  i[1819]);
assign l_40[1977]    = ( l_41 [3952] & !i[1819]) | ( l_41 [3953] &  i[1819]);
assign l_40[1978]    = ( l_41 [3954] & !i[1819]) | ( l_41 [3955] &  i[1819]);
assign l_40[1979]    = ( l_41 [3956] & !i[1819]) | ( l_41 [3957] &  i[1819]);
assign l_40[1980]    = ( l_41 [3958] & !i[1819]) | ( l_41 [3959] &  i[1819]);
assign l_40[1981]    = ( l_41 [3960] & !i[1819]) | ( l_41 [3961] &  i[1819]);
assign l_40[1982]    = ( l_41 [3962] & !i[1819]) | ( l_41 [3963] &  i[1819]);
assign l_40[1983]    = ( l_41 [3964] & !i[1819]) | ( l_41 [3965] &  i[1819]);
assign l_40[1984]    = ( l_41 [3966] & !i[1819]) | ( l_41 [3967] &  i[1819]);
assign l_40[1985]    = ( l_41 [3968] & !i[1819]) | ( l_41 [3969] &  i[1819]);
assign l_40[1986]    = ( l_41 [3970] & !i[1819]) | ( l_41 [3971] &  i[1819]);
assign l_40[1987]    = ( l_41 [3972] & !i[1819]) | ( l_41 [3973] &  i[1819]);
assign l_40[1988]    = ( l_41 [3974] & !i[1819]) | ( l_41 [3975] &  i[1819]);
assign l_40[1989]    = ( l_41 [3976] & !i[1819]) | ( l_41 [3977] &  i[1819]);
assign l_40[1990]    = ( l_41 [3978] & !i[1819]) | ( l_41 [3979] &  i[1819]);
assign l_40[1991]    = ( l_41 [3980] & !i[1819]) | ( l_41 [3981] &  i[1819]);
assign l_40[1992]    = ( l_41 [3982] & !i[1819]) | ( l_41 [3983] &  i[1819]);
assign l_40[1993]    = ( l_41 [3984] & !i[1819]) | ( l_41 [3985] &  i[1819]);
assign l_40[1994]    = ( l_41 [3986] & !i[1819]) | ( l_41 [3987] &  i[1819]);
assign l_40[1995]    = ( l_41 [3988] & !i[1819]) | ( l_41 [3989] &  i[1819]);
assign l_40[1996]    = ( l_41 [3990] & !i[1819]) | ( l_41 [3991] &  i[1819]);
assign l_40[1997]    = ( l_41 [3992] & !i[1819]) | ( l_41 [3993] &  i[1819]);
assign l_40[1998]    = ( l_41 [3994] & !i[1819]) | ( l_41 [3995] &  i[1819]);
assign l_40[1999]    = ( l_41 [3996] & !i[1819]) | ( l_41 [3997] &  i[1819]);
assign l_40[2000]    = ( l_41 [3998] & !i[1819]) | ( l_41 [3999] &  i[1819]);
assign l_40[2001]    = ( l_41 [4000] & !i[1819]) | ( l_41 [4001] &  i[1819]);
assign l_40[2002]    = ( l_41 [4002] & !i[1819]) | ( l_41 [4003] &  i[1819]);
assign l_40[2003]    = ( l_41 [4004] & !i[1819]) | ( l_41 [4005] &  i[1819]);
assign l_40[2004]    = ( l_41 [4006] & !i[1819]) | ( l_41 [4007] &  i[1819]);
assign l_40[2005]    = ( l_41 [4008] & !i[1819]) | ( l_41 [4009] &  i[1819]);
assign l_40[2006]    = ( l_41 [4010] & !i[1819]) | ( l_41 [4011] &  i[1819]);
assign l_40[2007]    = ( l_41 [4012] & !i[1819]) | ( l_41 [4013] &  i[1819]);
assign l_40[2008]    = ( l_41 [4014] & !i[1819]) | ( l_41 [4015] &  i[1819]);
assign l_40[2009]    = ( l_41 [4016] & !i[1819]) | ( l_41 [4017] &  i[1819]);
assign l_40[2010]    = ( l_41 [4018] & !i[1819]) | ( l_41 [4019] &  i[1819]);
assign l_40[2011]    = ( l_41 [4020] & !i[1819]) | ( l_41 [4021] &  i[1819]);
assign l_40[2012]    = ( l_41 [4022] & !i[1819]) | ( l_41 [4023] &  i[1819]);
assign l_40[2013]    = ( l_41 [4024] & !i[1819]) | ( l_41 [4025] &  i[1819]);
assign l_40[2014]    = ( l_41 [4026] & !i[1819]) | ( l_41 [4027] &  i[1819]);
assign l_40[2015]    = ( l_41 [4028] & !i[1819]) | ( l_41 [4029] &  i[1819]);
assign l_40[2016]    = ( l_41 [4030] & !i[1819]) | ( l_41 [4031] &  i[1819]);
assign l_40[2017]    = ( l_41 [4032] & !i[1819]) | ( l_41 [4033] &  i[1819]);
assign l_40[2018]    = ( l_41 [4034] & !i[1819]) | ( l_41 [4035] &  i[1819]);
assign l_40[2019]    = ( l_41 [4036] & !i[1819]) | ( l_41 [4037] &  i[1819]);
assign l_40[2020]    = ( l_41 [4038] & !i[1819]) | ( l_41 [4039] &  i[1819]);
assign l_40[2021]    = ( l_41 [4040] & !i[1819]) | ( l_41 [4041] &  i[1819]);
assign l_40[2022]    = ( l_41 [4042] & !i[1819]) | ( l_41 [4043] &  i[1819]);
assign l_40[2023]    = ( l_41 [4044] & !i[1819]) | ( l_41 [4045] &  i[1819]);
assign l_40[2024]    = ( l_41 [4046] & !i[1819]) | ( l_41 [4047] &  i[1819]);
assign l_40[2025]    = ( l_41 [4048] & !i[1819]) | ( l_41 [4049] &  i[1819]);
assign l_40[2026]    = ( l_41 [4050] & !i[1819]) | ( l_41 [4051] &  i[1819]);
assign l_40[2027]    = ( l_41 [4052] & !i[1819]) | ( l_41 [4053] &  i[1819]);
assign l_40[2028]    = ( l_41 [4054] & !i[1819]) | ( l_41 [4055] &  i[1819]);
assign l_40[2029]    = ( l_41 [4056] & !i[1819]) | ( l_41 [4057] &  i[1819]);
assign l_40[2030]    = ( l_41 [4058] & !i[1819]) | ( l_41 [4059] &  i[1819]);
assign l_40[2031]    = ( l_41 [4060] & !i[1819]) | ( l_41 [4061] &  i[1819]);
assign l_40[2032]    = ( l_41 [4062] & !i[1819]) | ( l_41 [4063] &  i[1819]);
assign l_40[2033]    = ( l_41 [4064] & !i[1819]) | ( l_41 [4065] &  i[1819]);
assign l_40[2034]    = ( l_41 [4066] & !i[1819]) | ( l_41 [4067] &  i[1819]);
assign l_40[2035]    = ( l_41 [4068] & !i[1819]) | ( l_41 [4069] &  i[1819]);
assign l_40[2036]    = ( l_41 [4070] & !i[1819]) | ( l_41 [4071] &  i[1819]);
assign l_40[2037]    = ( l_41 [4072] & !i[1819]) | ( l_41 [4073] &  i[1819]);
assign l_40[2038]    = ( l_41 [4074] & !i[1819]) | ( l_41 [4075] &  i[1819]);
assign l_40[2039]    = ( l_41 [4076] & !i[1819]) | ( l_41 [4077] &  i[1819]);
assign l_40[2040]    = ( l_41 [4078] & !i[1819]) | ( l_41 [4079] &  i[1819]);
assign l_40[2041]    = ( l_41 [4080] & !i[1819]) | ( l_41 [4081] &  i[1819]);
assign l_40[2042]    = ( l_41 [4082] & !i[1819]) | ( l_41 [4083] &  i[1819]);
assign l_40[2043]    = ( l_41 [4084] & !i[1819]) | ( l_41 [4085] &  i[1819]);
assign l_40[2044]    = ( l_41 [4086] & !i[1819]) | ( l_41 [4087] &  i[1819]);
assign l_40[2045]    = ( l_41 [4088] & !i[1819]) | ( l_41 [4089] &  i[1819]);
assign l_40[2046]    = ( l_41 [4090] & !i[1819]) | ( l_41 [4091] &  i[1819]);
assign l_40[2047]    = ( l_41 [4092] & !i[1819]) | ( l_41 [4093] &  i[1819]);
assign l_40[2048]    = ( l_41 [4094] & !i[1819]) | ( l_41 [4095] &  i[1819]);
assign l_40[2049]    = ( l_41 [4096] & !i[1819]) | ( l_41 [4097] &  i[1819]);
assign l_40[2050]    = ( l_41 [4098] & !i[1819]) | ( l_41 [4099] &  i[1819]);
assign l_40[2051]    = ( l_41 [4100] & !i[1819]) | ( l_41 [4101] &  i[1819]);
assign l_40[2052]    = ( l_41 [4102] & !i[1819]) | ( l_41 [4103] &  i[1819]);
assign l_40[2053]    = ( l_41 [4104] & !i[1819]) | ( l_41 [4105] &  i[1819]);
assign l_40[2054]    = ( l_41 [4106] & !i[1819]) | ( l_41 [4107] &  i[1819]);
assign l_40[2055]    = ( l_41 [4108] & !i[1819]) | ( l_41 [4109] &  i[1819]);
assign l_40[2056]    = ( l_41 [4110] & !i[1819]) | ( l_41 [4111] &  i[1819]);
assign l_40[2057]    = ( l_41 [4112] & !i[1819]) | ( l_41 [4113] &  i[1819]);
assign l_40[2058]    = ( l_41 [4114] & !i[1819]) | ( l_41 [4115] &  i[1819]);
assign l_40[2059]    = ( l_41 [4116] & !i[1819]) | ( l_41 [4117] &  i[1819]);
assign l_40[2060]    = ( l_41 [4118] & !i[1819]) | ( l_41 [4119] &  i[1819]);
assign l_40[2061]    = ( l_41 [4120] & !i[1819]) | ( l_41 [4121] &  i[1819]);
assign l_40[2062]    = ( l_41 [4122] & !i[1819]) | ( l_41 [4123] &  i[1819]);
assign l_40[2063]    = ( l_41 [4124] & !i[1819]) | ( l_41 [4125] &  i[1819]);
assign l_40[2064]    = ( l_41 [4126] & !i[1819]) | ( l_41 [4127] &  i[1819]);
assign l_40[2065]    = ( l_41 [4128] & !i[1819]) | ( l_41 [4129] &  i[1819]);
assign l_40[2066]    = ( l_41 [4130]);
assign l_40[2067]    = ( l_41 [4131]);
assign l_40[2068]    = ( l_41 [4132]);
assign l_40[2069]    = ( l_41 [4133]);
assign l_40[2070]    = ( l_41 [4134]);
assign l_40[2071]    = ( l_41 [4135]);
assign l_40[2072]    = ( l_41 [4136]);
assign l_40[2073]    = ( l_41 [4137]);
assign l_40[2074]    = ( l_41 [4138]);
assign l_40[2075]    = ( l_41 [4139]);
assign l_40[2076]    = ( l_41 [4140]);
assign l_40[2077]    = ( l_41 [4141]);
assign l_40[2078]    = ( l_41 [4142]);
assign l_40[2079]    = ( l_41 [4143]);
assign l_40[2080]    = ( l_41 [4144]);
assign l_40[2081]    = ( l_41 [4145]);
assign l_40[2082]    = ( l_41 [4146]);
assign l_40[2083]    = ( l_41 [4147]);
assign l_40[2084]    = ( l_41 [4148]);
assign l_40[2085]    = ( l_41 [4149]);
assign l_40[2086]    = ( l_41 [4150]);
assign l_40[2087]    = ( l_41 [4151]);
assign l_40[2088]    = ( l_41 [4152]);
assign l_40[2089]    = ( l_41 [4153]);
assign l_40[2090]    = ( l_41 [4154]);
assign l_40[2091]    = ( l_41 [4155]);
assign l_40[2092]    = ( l_41 [4156]);
assign l_40[2093]    = ( l_41 [4157]);
assign l_40[2094]    = ( l_41 [4158]);
assign l_40[2095]    = ( l_41 [4159]);
assign l_40[2096]    = ( l_41 [4160]);
assign l_40[2097]    = ( l_41 [4161]);
assign l_40[2098]    = ( l_41 [4162]);
assign l_40[2099]    = ( l_41 [4163]);
assign l_40[2100]    = ( l_41 [4164]);
assign l_40[2101]    = ( l_41 [4165]);
assign l_40[2102]    = ( l_41 [4166]);
assign l_40[2103]    = ( l_41 [4167]);
assign l_40[2104]    = ( l_41 [4168]);
assign l_40[2105]    = ( l_41 [4169]);
assign l_40[2106]    = ( l_41 [4170]);
assign l_40[2107]    = ( l_41 [4171]);
assign l_40[2108]    = ( l_41 [4172]);
assign l_40[2109]    = ( l_41 [4173]);
assign l_40[2110]    = ( l_41 [4174]);
assign l_40[2111]    = ( l_41 [4175]);
assign l_40[2112]    = ( l_41 [4176]);
assign l_40[2113]    = ( l_41 [4177]);
assign l_40[2114]    = ( l_41 [4178]);
assign l_40[2115]    = ( l_41 [4179]);
assign l_40[2116]    = ( l_41 [4180]);
assign l_40[2117]    = ( l_41 [4181]);
assign l_40[2118]    = ( l_41 [4182]);
assign l_40[2119]    = ( l_41 [4183]);
assign l_40[2120]    = ( l_41 [4184]);
assign l_40[2121]    = ( l_41 [4185]);
assign l_40[2122]    = ( l_41 [4186]);
assign l_40[2123]    = ( l_41 [4187]);
assign l_40[2124]    = ( l_41 [4188]);
assign l_40[2125]    = ( l_41 [4189]);
assign l_40[2126]    = ( l_41 [4190]);
assign l_40[2127]    = ( l_41 [4191]);
assign l_40[2128]    = ( l_41 [4192]);
assign l_40[2129]    = ( l_41 [4193]);
assign l_40[2130]    = ( l_41 [4194]);
assign l_40[2131]    = ( l_41 [4195]);
assign l_40[2132]    = ( l_41 [4196]);
assign l_40[2133]    = ( l_41 [4197]);
assign l_40[2134]    = ( l_41 [4198]);
assign l_40[2135]    = ( l_41 [4199]);
assign l_40[2136]    = ( l_41 [4200]);
assign l_40[2137]    = ( l_41 [4201]);
assign l_40[2138]    = ( l_41 [4202]);
assign l_40[2139]    = ( l_41 [4203]);
assign l_40[2140]    = ( l_41 [4204]);
assign l_40[2141]    = ( l_41 [4205]);
assign l_40[2142]    = ( l_41 [4206]);
assign l_40[2143]    = ( l_41 [4207]);
assign l_40[2144]    = ( l_41 [4208]);
assign l_40[2145]    = ( l_41 [4209]);
assign l_40[2146]    = ( l_41 [4210]);
assign l_40[2147]    = ( l_41 [4211]);
assign l_40[2148]    = ( l_41 [4212]);
assign l_40[2149]    = ( l_41 [4213]);
assign l_40[2150]    = ( l_41 [4214]);
assign l_40[2151]    = ( l_41 [4215]);
assign l_40[2152]    = ( l_41 [4216]);
assign l_40[2153]    = ( l_41 [4217]);
assign l_40[2154]    = ( l_41 [4218]);
assign l_40[2155]    = ( l_41 [4219]);
assign l_40[2156]    = ( l_41 [4220]);
assign l_40[2157]    = ( l_41 [4221]);
assign l_40[2158]    = ( l_41 [4222]);
assign l_40[2159]    = ( l_41 [4223]);
assign l_40[2160]    = ( l_41 [4224]);
assign l_40[2161]    = ( l_41 [4225]);
assign l_40[2162]    = ( l_41 [4226]);
assign l_40[2163]    = ( l_41 [4227]);
assign l_40[2164]    = ( l_41 [4228]);
assign l_40[2165]    = ( l_41 [4229]);
assign l_40[2166]    = ( l_41 [4230]);
assign l_40[2167]    = ( l_41 [4231]);
assign l_40[2168]    = ( l_41 [4232]);
assign l_40[2169]    = ( l_41 [4233]);
assign l_40[2170]    = ( l_41 [4234]);
assign l_40[2171]    = ( l_41 [4235]);
assign l_40[2172]    = ( l_41 [4236]);
assign l_40[2173]    = ( l_41 [4237]);
assign l_40[2174]    = ( l_41 [4238]);
assign l_40[2175]    = ( l_41 [4239]);
assign l_40[2176]    = ( l_41 [4240]);
assign l_40[2177]    = ( l_41 [4241]);
assign l_40[2178]    = ( l_41 [4242]);
assign l_40[2179]    = ( l_41 [4243]);
assign l_40[2180]    = ( l_41 [4244]);
assign l_40[2181]    = ( l_41 [4245]);
assign l_40[2182]    = ( l_41 [4246]);
assign l_40[2183]    = ( l_41 [4247]);
assign l_40[2184]    = ( l_41 [4248]);
assign l_40[2185]    = ( l_41 [4249]);
assign l_40[2186]    = ( l_41 [4250]);
assign l_40[2187]    = ( l_41 [4251]);
assign l_40[2188]    = ( l_41 [4252]);
assign l_40[2189]    = ( l_41 [4253]);
assign l_40[2190]    = ( l_41 [4254]);
assign l_40[2191]    = ( l_41 [4255]);
assign l_40[2192]    = ( l_41 [4256]);
assign l_40[2193]    = ( l_41 [4257]);
assign l_40[2194]    = ( l_41 [4258]);
assign l_40[2195]    = ( l_41 [4259]);
assign l_40[2196]    = ( l_41 [4260]);
assign l_40[2197]    = ( l_41 [4261]);
assign l_40[2198]    = ( l_41 [4262]);
assign l_40[2199]    = ( l_41 [4263]);
assign l_40[2200]    = ( l_41 [4264]);
assign l_40[2201]    = ( l_41 [4265]);
assign l_40[2202]    = ( l_41 [4266]);
assign l_40[2203]    = ( l_41 [4267]);
assign l_40[2204]    = ( l_41 [4268]);
assign l_40[2205]    = ( l_41 [4269]);
assign l_40[2206]    = ( l_41 [4270]);
assign l_40[2207]    = ( l_41 [4271]);
assign l_40[2208]    = ( l_41 [4272]);
assign l_40[2209]    = ( l_41 [4273]);
assign l_40[2210]    = ( l_41 [4274]);
assign l_40[2211]    = ( l_41 [4275]);
assign l_40[2212]    = ( l_41 [4276]);
assign l_40[2213]    = ( l_41 [4277]);
assign l_40[2214]    = ( l_41 [4278]);
assign l_40[2215]    = ( l_41 [4279]);
assign l_40[2216]    = ( l_41 [4280]);
assign l_40[2217]    = ( l_41 [4281]);
assign l_40[2218]    = ( l_41 [4282]);
assign l_40[2219]    = ( l_41 [4283]);
assign l_40[2220]    = ( l_41 [4284]);
assign l_40[2221]    = ( l_41 [4285]);
assign l_40[2222]    = ( l_41 [4286]);
assign l_40[2223]    = ( l_41 [4287]);
assign l_40[2224]    = ( l_41 [4288]);
assign l_40[2225]    = ( l_41 [4289]);
assign l_40[2226]    = ( l_41 [4290]);
assign l_40[2227]    = ( l_41 [4291]);
assign l_40[2228]    = ( l_41 [4292]);
assign l_40[2229]    = ( l_41 [4293]);
assign l_40[2230]    = ( l_41 [4294]);
assign l_40[2231]    = ( l_41 [4295]);
assign l_40[2232]    = ( l_41 [4296]);
assign l_40[2233]    = ( l_41 [4297]);
assign l_40[2234]    = ( l_41 [4298]);
assign l_40[2235]    = ( l_41 [4299]);
assign l_40[2236]    = ( l_41 [4300]);
assign l_40[2237]    = ( l_41 [4301]);
assign l_40[2238]    = ( l_41 [4302]);
assign l_40[2239]    = ( l_41 [4303]);
assign l_40[2240]    = ( l_41 [4304]);
assign l_40[2241]    = ( l_41 [4305]);
assign l_40[2242]    = ( l_41 [4306]);
assign l_40[2243]    = ( l_41 [4307]);
assign l_40[2244]    = ( l_41 [4308]);
assign l_40[2245]    = ( l_41 [4309]);
assign l_40[2246]    = ( l_41 [4310]);
assign l_40[2247]    = ( l_41 [4311]);
assign l_40[2248]    = ( l_41 [4312]);
assign l_40[2249]    = ( l_41 [4313]);
assign l_40[2250]    = ( l_41 [4314]);
assign l_40[2251]    = ( l_41 [4315]);
assign l_40[2252]    = ( l_41 [4316]);
assign l_40[2253]    = ( l_41 [4317]);
assign l_40[2254]    = ( l_41 [4318]);
assign l_40[2255]    = ( l_41 [4319]);
assign l_40[2256]    = ( l_41 [4320]);
assign l_40[2257]    = ( l_41 [4321]);
assign l_40[2258]    = ( l_41 [4322]);
assign l_40[2259]    = ( l_41 [4323]);
assign l_40[2260]    = ( l_41 [4324]);
assign l_40[2261]    = ( l_41 [4325]);
assign l_40[2262]    = ( l_41 [4326]);
assign l_40[2263]    = ( l_41 [4327]);
assign l_40[2264]    = ( l_41 [4328]);
assign l_40[2265]    = ( l_41 [4329]);
assign l_40[2266]    = ( l_41 [4330]);
assign l_40[2267]    = ( l_41 [4331]);
assign l_40[2268]    = ( l_41 [4332]);
assign l_40[2269]    = ( l_41 [4333]);
assign l_40[2270]    = ( l_41 [4334]);
assign l_40[2271]    = ( l_41 [4335]);
assign l_40[2272]    = ( l_41 [4336]);
assign l_40[2273]    = ( l_41 [4337]);
assign l_40[2274]    = ( l_41 [4338]);
assign l_40[2275]    = ( l_41 [4339]);
assign l_40[2276]    = ( l_41 [4340]);
assign l_40[2277]    = ( l_41 [4341]);
assign l_40[2278]    = ( l_41 [4342]);
assign l_40[2279]    = ( l_41 [4343]);
assign l_40[2280]    = ( l_41 [4344]);
assign l_40[2281]    = ( l_41 [4345]);
assign l_40[2282]    = ( l_41 [4346]);
assign l_40[2283]    = ( l_41 [4347]);
assign l_40[2284]    = ( l_41 [4348]);
assign l_40[2285]    = ( l_41 [4349]);
assign l_40[2286]    = ( l_41 [4350]);
assign l_40[2287]    = ( l_41 [4351]);
assign l_40[2288]    = ( l_41 [4352]);
assign l_40[2289]    = ( l_41 [4353]);
assign l_40[2290]    = ( l_41 [4354]);
assign l_40[2291]    = ( l_41 [4355]);
assign l_40[2292]    = ( l_41 [4356]);
assign l_40[2293]    = ( l_41 [4357]);
assign l_40[2294]    = ( l_41 [4358]);
assign l_40[2295]    = ( l_41 [4359]);
assign l_40[2296]    = ( l_41 [4360]);
assign l_40[2297]    = ( l_41 [4361]);
assign l_40[2298]    = ( l_41 [4362]);
assign l_40[2299]    = ( l_41 [4363]);
assign l_40[2300]    = ( l_41 [4364]);
assign l_40[2301]    = ( l_41 [4365]);
assign l_40[2302]    = ( l_41 [4366]);
assign l_40[2303]    = ( l_41 [4367]);
assign l_40[2304]    = ( l_41 [4368]);
assign l_40[2305]    = ( l_41 [4369]);
assign l_40[2306]    = ( l_41 [4370]);
assign l_40[2307]    = ( l_41 [4371]);
assign l_40[2308]    = ( l_41 [4372]);
assign l_40[2309]    = ( l_41 [4373]);
assign l_40[2310]    = ( l_41 [4374]);
assign l_40[2311]    = ( l_41 [4375]);
assign l_40[2312]    = ( l_41 [4376]);
assign l_40[2313]    = ( l_41 [4377]);
assign l_40[2314]    = ( l_41 [4378]);
assign l_40[2315]    = ( l_41 [4379]);
assign l_40[2316]    = ( l_41 [4380]);
assign l_40[2317]    = ( l_41 [4381]);
assign l_40[2318]    = ( l_41 [4382]);
assign l_40[2319]    = ( l_41 [4383]);
assign l_40[2320]    = ( l_41 [4384]);
assign l_40[2321]    = ( l_41 [4385]);
assign l_40[2322]    = ( l_41 [4386]);
assign l_40[2323]    = ( l_41 [4387]);
assign l_40[2324]    = ( l_41 [4388]);
assign l_40[2325]    = ( l_41 [4389]);
assign l_40[2326]    = ( l_41 [4390]);
assign l_40[2327]    = ( l_41 [4391]);
assign l_40[2328]    = ( l_41 [4392]);
assign l_40[2329]    = ( l_41 [4393]);
assign l_40[2330]    = ( l_41 [4394]);
assign l_40[2331]    = ( l_41 [4395]);
assign l_40[2332]    = ( l_41 [4396]);
assign l_40[2333]    = ( l_41 [4397]);
assign l_40[2334]    = ( l_41 [4398]);
assign l_40[2335]    = ( l_41 [4399]);
assign l_40[2336]    = ( l_41 [4400]);
assign l_40[2337]    = ( l_41 [4401]);
assign l_40[2338]    = ( l_41 [4402]);
assign l_40[2339]    = ( l_41 [4403]);
assign l_40[2340]    = ( l_41 [4404]);
assign l_40[2341]    = ( l_41 [4405]);
assign l_40[2342]    = ( l_41 [4406]);
assign l_40[2343]    = ( l_41 [4407]);
assign l_40[2344]    = ( l_41 [4408]);
assign l_40[2345]    = ( l_41 [4409]);
assign l_40[2346]    = ( l_41 [4410]);
assign l_40[2347]    = ( l_41 [4411]);
assign l_40[2348]    = ( l_41 [4412]);
assign l_40[2349]    = ( l_41 [4413]);
assign l_40[2350]    = ( l_41 [4414]);
assign l_40[2351]    = ( l_41 [4415]);
assign l_40[2352]    = ( l_41 [4416]);
assign l_40[2353]    = ( l_41 [4417]);
assign l_40[2354]    = ( l_41 [4418]);
assign l_40[2355]    = ( l_41 [4419]);
assign l_40[2356]    = ( l_41 [4420]);
assign l_40[2357]    = ( l_41 [4421]);
assign l_40[2358]    = ( l_41 [4422]);
assign l_40[2359]    = ( l_41 [4423]);
assign l_40[2360]    = ( l_41 [4424]);
assign l_40[2361]    = ( l_41 [4425]);
assign l_40[2362]    = ( l_41 [4426]);
assign l_40[2363]    = ( l_41 [4427]);
assign l_40[2364]    = ( l_41 [4428]);
assign l_40[2365]    = ( l_41 [4429]);
assign l_40[2366]    = ( l_41 [4430]);
assign l_40[2367]    = ( l_41 [4431]);
assign l_40[2368]    = ( l_41 [4432]);
assign l_40[2369]    = ( l_41 [4433]);
assign l_40[2370]    = ( l_41 [4434]);
assign l_40[2371]    = ( l_41 [4435]);
assign l_40[2372]    = ( l_41 [4436]);
assign l_40[2373]    = ( l_41 [4437]);
assign l_40[2374]    = ( l_41 [4438]);
assign l_40[2375]    = ( l_41 [4439]);
assign l_40[2376]    = ( l_41 [4440]);
assign l_40[2377]    = ( l_41 [4441]);
assign l_40[2378]    = ( l_41 [4442]);
assign l_40[2379]    = ( l_41 [4443]);
assign l_40[2380]    = ( l_41 [4444]);
assign l_40[2381]    = ( l_41 [4445]);
assign l_40[2382]    = ( l_41 [4446]);
assign l_40[2383]    = ( l_41 [4447]);
assign l_40[2384]    = ( l_41 [4448]);
assign l_40[2385]    = ( l_41 [4449]);
assign l_40[2386]    = ( l_41 [4450]);
assign l_40[2387]    = ( l_41 [4451]);
assign l_40[2388]    = ( l_41 [4452]);
assign l_40[2389]    = ( l_41 [4453]);
assign l_40[2390]    = ( l_41 [4454]);
assign l_40[2391]    = ( l_41 [4455]);
assign l_40[2392]    = ( l_41 [4456]);
assign l_40[2393]    = ( l_41 [4457]);
assign l_40[2394]    = ( l_41 [4458]);
assign l_40[2395]    = ( l_41 [4459]);
assign l_40[2396]    = ( l_41 [4460]);
assign l_40[2397]    = ( l_41 [4461]);
assign l_40[2398]    = ( l_41 [4462]);
assign l_40[2399]    = ( l_41 [4463]);
assign l_40[2400]    = ( l_41 [4464]);
assign l_40[2401]    = ( l_41 [4465]);
assign l_40[2402]    = ( l_41 [4466]);
assign l_40[2403]    = ( l_41 [4467]);
assign l_40[2404]    = ( l_41 [4468]);
assign l_40[2405]    = ( l_41 [4469]);
assign l_40[2406]    = ( l_41 [4470]);
assign l_40[2407]    = ( l_41 [4471]);
assign l_40[2408]    = ( l_41 [4472]);
assign l_40[2409]    = ( l_41 [4473]);
assign l_40[2410]    = ( l_41 [4474]);
assign l_40[2411]    = ( l_41 [4475]);
assign l_40[2412]    = ( l_41 [4476]);
assign l_40[2413]    = ( l_41 [4477]);
assign l_40[2414]    = ( l_41 [4478]);
assign l_40[2415]    = ( l_41 [4479]);
assign l_40[2416]    = ( l_41 [4480]);
assign l_40[2417]    = ( l_41 [4481]);
assign l_40[2418]    = ( l_41 [4482]);
assign l_40[2419]    = ( l_41 [4483]);
assign l_40[2420]    = ( l_41 [4484]);
assign l_40[2421]    = ( l_41 [4485]);
assign l_40[2422]    = ( l_41 [4486]);
assign l_40[2423]    = ( l_41 [4487]);
assign l_40[2424]    = ( l_41 [4488]);
assign l_40[2425]    = ( l_41 [4489]);
assign l_40[2426]    = ( l_41 [4490]);
assign l_40[2427]    = ( l_41 [4491]);
assign l_40[2428]    = ( l_41 [4492]);
assign l_40[2429]    = ( l_41 [4493]);
assign l_40[2430]    = ( l_41 [4494]);
assign l_40[2431]    = ( l_41 [4495]);
assign l_40[2432]    = ( l_41 [4496]);
assign l_40[2433]    = ( l_41 [4497]);
assign l_40[2434]    = ( l_41 [4498]);
assign l_40[2435]    = ( l_41 [4499]);
assign l_40[2436]    = ( l_41 [4500]);
assign l_40[2437]    = ( l_41 [4501]);
assign l_40[2438]    = ( l_41 [4502]);
assign l_40[2439]    = ( l_41 [4503]);
assign l_40[2440]    = ( l_41 [4504]);
assign l_40[2441]    = ( l_41 [4505]);
assign l_40[2442]    = ( l_41 [4506]);
assign l_40[2443]    = ( l_41 [4507]);
assign l_40[2444]    = ( l_41 [4508]);
assign l_40[2445]    = ( l_41 [4509]);
assign l_40[2446]    = ( l_41 [4510]);
assign l_40[2447]    = ( l_41 [4511]);
assign l_40[2448]    = ( l_41 [4512]);
assign l_40[2449]    = ( l_41 [4513]);
assign l_40[2450]    = ( l_41 [4514]);
assign l_40[2451]    = ( l_41 [4515]);
assign l_40[2452]    = ( l_41 [4516]);
assign l_40[2453]    = ( l_41 [4517]);
assign l_40[2454]    = ( l_41 [4518]);
assign l_40[2455]    = ( l_41 [4519]);
assign l_40[2456]    = ( l_41 [4520]);
assign l_40[2457]    = ( l_41 [4521]);
assign l_40[2458]    = ( l_41 [4522]);
assign l_40[2459]    = ( l_41 [4523]);
assign l_40[2460]    = ( l_41 [4524]);
assign l_40[2461]    = ( l_41 [4525]);
assign l_40[2462]    = ( l_41 [4526]);
assign l_40[2463]    = ( l_41 [4527]);
assign l_40[2464]    = ( l_41 [4528]);
assign l_40[2465]    = ( l_41 [4529]);
assign l_40[2466]    = ( l_41 [4530]);
assign l_40[2467]    = ( l_41 [4531]);
assign l_40[2468]    = ( l_41 [4532]);
assign l_40[2469]    = ( l_41 [4533]);
assign l_40[2470]    = ( l_41 [4534]);
assign l_40[2471]    = ( l_41 [4535]);
assign l_40[2472]    = ( l_41 [4536]);
assign l_40[2473]    = ( l_41 [4537]);
assign l_40[2474]    = ( l_41 [4538]);
assign l_40[2475]    = ( l_41 [4539]);
assign l_40[2476]    = ( l_41 [4540]);
assign l_40[2477]    = ( l_41 [4541]);
assign l_40[2478]    = ( l_41 [4542]);
assign l_40[2479]    = ( l_41 [4543]);
assign l_40[2480]    = ( l_41 [4544]);
assign l_40[2481]    = ( l_41 [4545]);
assign l_40[2482]    = ( l_41 [4546]);
assign l_40[2483]    = ( l_41 [4547]);
assign l_40[2484]    = ( l_41 [4548]);
assign l_40[2485]    = ( l_41 [4549]);
assign l_40[2486]    = ( l_41 [4550]);
assign l_40[2487]    = ( l_41 [4551]);
assign l_40[2488]    = ( l_41 [4552]);
assign l_40[2489]    = ( l_41 [4553]);
assign l_40[2490]    = ( l_41 [4554]);
assign l_40[2491]    = ( l_41 [4555]);
assign l_40[2492]    = ( l_41 [4556]);
assign l_40[2493]    = ( l_41 [4557]);
assign l_40[2494]    = ( l_41 [4558]);
assign l_40[2495]    = ( l_41 [4559]);
assign l_40[2496]    = ( l_41 [4560]);
assign l_40[2497]    = ( l_41 [4561]);
assign l_40[2498]    = ( l_41 [4562]);
assign l_40[2499]    = ( l_41 [4563]);
assign l_40[2500]    = ( l_41 [4564]);
assign l_40[2501]    = ( l_41 [4565]);
assign l_40[2502]    = ( l_41 [4566]);
assign l_40[2503]    = ( l_41 [4567]);
assign l_40[2504]    = ( l_41 [4568]);
assign l_40[2505]    = ( l_41 [4569]);
assign l_40[2506]    = ( l_41 [4570]);
assign l_40[2507]    = ( l_41 [4571]);
assign l_40[2508]    = ( l_41 [4572]);
assign l_40[2509]    = ( l_41 [4573]);
assign l_40[2510]    = ( l_41 [4574]);
assign l_40[2511]    = ( l_41 [4575]);
assign l_40[2512]    = ( l_41 [4576]);
assign l_40[2513]    = ( l_41 [4577]);
assign l_40[2514]    = ( l_41 [4578]);
assign l_40[2515]    = ( l_41 [4579]);
assign l_40[2516]    = ( l_41 [4580]);
assign l_40[2517]    = ( l_41 [4581]);
assign l_40[2518]    = ( l_41 [4582]);
assign l_40[2519]    = ( l_41 [4583]);
assign l_40[2520]    = ( l_41 [4584]);
assign l_40[2521]    = ( l_41 [4585]);
assign l_40[2522]    = ( l_41 [4586]);
assign l_40[2523]    = ( l_41 [4587]);
assign l_40[2524]    = ( l_41 [4588]);
assign l_40[2525]    = ( l_41 [4589]);
assign l_40[2526]    = ( l_41 [4590]);
assign l_40[2527]    = ( l_41 [4591]);
assign l_40[2528]    = ( l_41 [4592]);
assign l_40[2529]    = ( l_41 [4593]);
assign l_40[2530]    = ( l_41 [4594]);
assign l_40[2531]    = ( l_41 [4595]);
assign l_40[2532]    = ( l_41 [4596]);
assign l_40[2533]    = ( l_41 [4597]);
assign l_40[2534]    = ( l_41 [4598]);
assign l_40[2535]    = ( l_41 [4599]);
assign l_40[2536]    = ( l_41 [4600]);
assign l_40[2537]    = ( l_41 [4601]);
assign l_40[2538]    = ( l_41 [4602]);
assign l_40[2539]    = ( l_41 [4603]);
assign l_40[2540]    = ( l_41 [4604]);
assign l_40[2541]    = ( l_41 [4605]);
assign l_40[2542]    = ( l_41 [4606]);
assign l_40[2543]    = ( l_41 [4607]);
assign l_40[2544]    = ( l_41 [4608]);
assign l_40[2545]    = ( l_41 [4609]);
assign l_40[2546]    = ( l_41 [4610]);
assign l_40[2547]    = ( l_41 [4611]);
assign l_40[2548]    = ( l_41 [4612]);
assign l_40[2549]    = ( l_41 [4613]);
assign l_40[2550]    = ( l_41 [4614]);
assign l_40[2551]    = ( l_41 [4615]);
assign l_40[2552]    = ( l_41 [4616]);
assign l_40[2553]    = ( l_41 [4617]);
assign l_40[2554]    = ( l_41 [4618]);
assign l_40[2555]    = ( l_41 [4619]);
assign l_40[2556]    = ( l_41 [4620]);
assign l_40[2557]    = ( l_41 [4621]);
assign l_40[2558]    = ( l_41 [4622]);
assign l_40[2559]    = ( l_41 [4623]);
assign l_40[2560]    = ( l_41 [4624]);
assign l_40[2561]    = ( l_41 [4625]);
assign l_40[2562]    = ( l_41 [4626]);
assign l_40[2563]    = ( l_41 [4627]);
assign l_40[2564]    = ( l_41 [4628]);
assign l_40[2565]    = ( l_41 [4629]);
assign l_40[2566]    = ( l_41 [4630]);
assign l_40[2567]    = ( l_41 [4631]);
assign l_40[2568]    = ( l_41 [4632]);
assign l_40[2569]    = ( l_41 [4633]);
assign l_40[2570]    = ( l_41 [4634]);
assign l_40[2571]    = ( l_41 [4635]);
assign l_40[2572]    = ( l_41 [4636]);
assign l_40[2573]    = ( l_41 [4637]);
assign l_40[2574]    = ( l_41 [4638]);
assign l_40[2575]    = ( l_41 [4639]);
assign l_40[2576]    = ( l_41 [4640]);
assign l_40[2577]    = ( l_41 [4641]);
assign l_40[2578]    = ( l_41 [4642]);
assign l_40[2579]    = ( l_41 [4643]);
assign l_40[2580]    = ( l_41 [4644]);
assign l_40[2581]    = ( l_41 [4645]);
assign l_40[2582]    = ( l_41 [4646]);
assign l_40[2583]    = ( l_41 [4647]);
assign l_40[2584]    = ( l_41 [4648]);
assign l_40[2585]    = ( l_41 [4649]);
assign l_40[2586]    = ( l_41 [4650]);
assign l_40[2587]    = ( l_41 [4651]);
assign l_40[2588]    = ( l_41 [4652]);
assign l_40[2589]    = ( l_41 [4653]);
assign l_40[2590]    = ( l_41 [4654]);
assign l_40[2591]    = ( l_41 [4655]);
assign l_40[2592]    = ( l_41 [4656]);
assign l_40[2593]    = ( l_41 [4657]);
assign l_40[2594]    = ( l_41 [4658]);
assign l_40[2595]    = ( l_41 [4659]);
assign l_40[2596]    = ( l_41 [4660]);
assign l_40[2597]    = ( l_41 [4661]);
assign l_40[2598]    = ( l_41 [4662]);
assign l_40[2599]    = ( l_41 [4663]);
assign l_40[2600]    = ( l_41 [4664]);
assign l_40[2601]    = ( l_41 [4665]);
assign l_40[2602]    = ( l_41 [4666]);
assign l_40[2603]    = ( l_41 [4667]);
assign l_40[2604]    = ( l_41 [4668]);
assign l_40[2605]    = ( l_41 [4669]);
assign l_40[2606]    = ( l_41 [4670]);
assign l_40[2607]    = ( l_41 [4671]);
assign l_40[2608]    = ( l_41 [4672]);
assign l_40[2609]    = ( l_41 [4673]);
assign l_40[2610]    = ( l_41 [4674]);
assign l_40[2611]    = ( l_41 [4675]);
assign l_40[2612]    = ( l_41 [4676]);
assign l_40[2613]    = ( l_41 [4677]);
assign l_40[2614]    = ( l_41 [4678]);
assign l_40[2615]    = ( l_41 [4679]);
assign l_40[2616]    = ( l_41 [4680]);
assign l_40[2617]    = ( l_41 [4681]);
assign l_40[2618]    = ( l_41 [4682]);
assign l_40[2619]    = ( l_41 [4683]);
assign l_40[2620]    = ( l_41 [4684]);
assign l_40[2621]    = ( l_41 [4685]);
assign l_40[2622]    = ( l_41 [4686]);
assign l_40[2623]    = ( l_41 [4687]);
assign l_40[2624]    = ( l_41 [4688]);
assign l_40[2625]    = ( l_41 [4689]);
assign l_40[2626]    = ( l_41 [4690]);
assign l_40[2627]    = ( l_41 [4691]);
assign l_40[2628]    = ( l_41 [4692]);
assign l_40[2629]    = ( l_41 [4693]);
assign l_40[2630]    = ( l_41 [4694]);
assign l_40[2631]    = ( l_41 [4695]);
assign l_40[2632]    = ( l_41 [4696]);
assign l_40[2633]    = ( l_41 [4697]);
assign l_40[2634]    = ( l_41 [4698]);
assign l_40[2635]    = ( l_41 [4699]);
assign l_40[2636]    = ( l_41 [4700]);
assign l_40[2637]    = ( l_41 [4701]);
assign l_40[2638]    = ( l_41 [4702]);
assign l_40[2639]    = ( l_41 [4703]);
assign l_40[2640]    = ( l_41 [4704]);
assign l_40[2641]    = ( l_41 [4705]);
assign l_40[2642]    = ( l_41 [4706]);
assign l_40[2643]    = ( l_41 [4707]);
assign l_40[2644]    = ( l_41 [4708]);
assign l_40[2645]    = ( l_41 [4709]);
assign l_40[2646]    = ( l_41 [4710]);
assign l_40[2647]    = ( l_41 [4711]);
assign l_40[2648]    = ( l_41 [4712]);
assign l_40[2649]    = ( l_41 [4713]);
assign l_40[2650]    = ( l_41 [4714]);
assign l_40[2651]    = ( l_41 [4715]);
assign l_40[2652]    = ( l_41 [4716]);
assign l_40[2653]    = ( l_41 [4717]);
assign l_40[2654]    = ( l_41 [4718]);
assign l_40[2655]    = ( l_41 [4719]);
assign l_40[2656]    = ( l_41 [4720]);
assign l_40[2657]    = ( l_41 [4721]);
assign l_40[2658]    = ( l_41 [4722]);
assign l_40[2659]    = ( l_41 [4723]);
assign l_40[2660]    = ( l_41 [4724]);
assign l_40[2661]    = ( l_41 [4725]);
assign l_40[2662]    = ( l_41 [4726]);
assign l_40[2663]    = ( l_41 [4727]);
assign l_40[2664]    = ( l_41 [4728]);
assign l_40[2665]    = ( l_41 [4729]);
assign l_40[2666]    = ( l_41 [4730]);
assign l_40[2667]    = ( l_41 [4731]);
assign l_40[2668]    = ( l_41 [4732]);
assign l_40[2669]    = ( l_41 [4733]);
assign l_40[2670]    = ( l_41 [4734]);
assign l_40[2671]    = ( l_41 [4735]);
assign l_40[2672]    = ( l_41 [4736]);
assign l_40[2673]    = ( l_41 [4737]);
assign l_40[2674]    = ( l_41 [4738]);
assign l_40[2675]    = ( l_41 [4739]);
assign l_40[2676]    = ( l_41 [4740]);
assign l_40[2677]    = ( l_41 [4741]);
assign l_40[2678]    = ( l_41 [4742]);
assign l_40[2679]    = ( l_41 [4743]);
assign l_40[2680]    = ( l_41 [4744]);
assign l_40[2681]    = ( l_41 [4745]);
assign l_40[2682]    = ( l_41 [4746]);
assign l_40[2683]    = ( l_41 [4747]);
assign l_40[2684]    = ( l_41 [4748]);
assign l_40[2685]    = ( l_41 [4749]);
assign l_40[2686]    = ( l_41 [4750]);
assign l_40[2687]    = ( l_41 [4751]);
assign l_40[2688]    = ( l_41 [4752]);
assign l_40[2689]    = ( l_41 [4753]);
assign l_40[2690]    = ( l_41 [4754]);
assign l_40[2691]    = ( l_41 [4755]);
assign l_40[2692]    = ( l_41 [4756]);
assign l_40[2693]    = ( l_41 [4757]);
assign l_40[2694]    = ( l_41 [4758]);
assign l_40[2695]    = ( l_41 [4759]);
assign l_40[2696]    = ( l_41 [4760]);
assign l_40[2697]    = ( l_41 [4761]);
assign l_40[2698]    = ( l_41 [4762]);
assign l_40[2699]    = ( l_41 [4763]);
assign l_40[2700]    = ( l_41 [4764]);
assign l_40[2701]    = ( l_41 [4765]);
assign l_40[2702]    = ( l_41 [4766]);
assign l_40[2703]    = ( l_41 [4767]);
assign l_40[2704]    = ( l_41 [4768]);
assign l_40[2705]    = ( l_41 [4769]);
assign l_40[2706]    = ( l_41 [4770]);
assign l_40[2707]    = ( l_41 [4771]);
assign l_40[2708]    = ( l_41 [4772]);
assign l_40[2709]    = ( l_41 [4773]);
assign l_40[2710]    = ( l_41 [4774]);
assign l_40[2711]    = ( l_41 [4775]);
assign l_40[2712]    = ( l_41 [4776]);
assign l_40[2713]    = ( l_41 [4777]);
assign l_40[2714]    = ( l_41 [4778]);
assign l_40[2715]    = ( l_41 [4779]);
assign l_40[2716]    = ( l_41 [4780]);
assign l_40[2717]    = ( l_41 [4781]);
assign l_40[2718]    = ( l_41 [4782]);
assign l_40[2719]    = ( l_41 [4783]);
assign l_40[2720]    = ( l_41 [4784]);
assign l_40[2721]    = ( l_41 [4785]);
assign l_40[2722]    = ( l_41 [4786]);
assign l_40[2723]    = ( l_41 [4787]);
assign l_40[2724]    = ( l_41 [4788]);
assign l_40[2725]    = ( l_41 [4789]);
assign l_40[2726]    = ( l_41 [4790]);
assign l_40[2727]    = ( l_41 [4791]);
assign l_40[2728]    = ( l_41 [4792]);
assign l_40[2729]    = ( l_41 [4793]);
assign l_40[2730]    = ( l_41 [4794]);
assign l_40[2731]    = ( l_41 [4795]);
assign l_40[2732]    = ( l_41 [4796]);
assign l_40[2733]    = ( l_41 [4797]);
assign l_40[2734]    = ( l_41 [4798]);
assign l_40[2735]    = ( l_41 [4799]);
assign l_40[2736]    = ( l_41 [4800]);
assign l_40[2737]    = ( l_41 [4801]);
assign l_40[2738]    = ( l_41 [4802]);
assign l_40[2739]    = ( l_41 [4803]);
assign l_40[2740]    = ( l_41 [4804]);
assign l_40[2741]    = ( l_41 [4805]);
assign l_40[2742]    = ( l_41 [4806]);
assign l_40[2743]    = ( l_41 [4807]);
assign l_40[2744]    = ( l_41 [4808]);
assign l_40[2745]    = ( l_41 [4809]);
assign l_40[2746]    = ( l_41 [4810]);
assign l_40[2747]    = ( l_41 [4811]);
assign l_40[2748]    = ( l_41 [4812]);
assign l_40[2749]    = ( l_41 [4813]);
assign l_40[2750]    = ( l_41 [4814]);
assign l_40[2751]    = ( l_41 [4815]);
assign l_40[2752]    = ( l_41 [4816]);
assign l_40[2753]    = ( l_41 [4817]);
assign l_40[2754]    = ( l_41 [4818]);
assign l_40[2755]    = ( l_41 [4819]);
assign l_40[2756]    = ( l_41 [4820]);
assign l_40[2757]    = ( l_41 [4821]);
assign l_40[2758]    = ( l_41 [4822]);
assign l_40[2759]    = ( l_41 [4823]);
assign l_40[2760]    = ( l_41 [4824]);
assign l_40[2761]    = ( l_41 [4825]);
assign l_40[2762]    = ( l_41 [4826]);
assign l_40[2763]    = ( l_41 [4827]);
assign l_40[2764]    = ( l_41 [4828]);
assign l_40[2765]    = ( l_41 [4829]);
assign l_40[2766]    = ( l_41 [4830]);
assign l_40[2767]    = ( l_41 [4831]);
assign l_40[2768]    = ( l_41 [4832]);
assign l_40[2769]    = ( l_41 [4833]);
assign l_40[2770]    = ( l_41 [4834]);
assign l_40[2771]    = ( l_41 [4835]);
assign l_40[2772]    = ( l_41 [4836]);
assign l_40[2773]    = ( l_41 [4837]);
assign l_40[2774]    = ( l_41 [4838]);
assign l_40[2775]    = ( l_41 [4839]);
assign l_40[2776]    = ( l_41 [4840]);
assign l_40[2777]    = ( l_41 [4841]);
assign l_40[2778]    = ( l_41 [4842]);
assign l_40[2779]    = ( l_41 [4843]);
assign l_40[2780]    = ( l_41 [4844]);
assign l_40[2781]    = ( l_41 [4845]);
assign l_40[2782]    = ( l_41 [4846]);
assign l_40[2783]    = ( l_41 [4847]);
assign l_40[2784]    = ( l_41 [4848]);
assign l_40[2785]    = ( l_41 [4849]);
assign l_40[2786]    = ( l_41 [4850]);
assign l_40[2787]    = ( l_41 [4851]);
assign l_40[2788]    = ( l_41 [4852]);
assign l_40[2789]    = ( l_41 [4853]);
assign l_40[2790]    = ( l_41 [4854]);
assign l_40[2791]    = ( l_41 [4855]);
assign l_40[2792]    = ( l_41 [4856]);
assign l_40[2793]    = ( l_41 [4857]);
assign l_40[2794]    = ( l_41 [4858]);
assign l_40[2795]    = ( l_41 [4859]);
assign l_40[2796]    = ( l_41 [4860]);
assign l_40[2797]    = ( l_41 [4861]);
assign l_40[2798]    = ( l_41 [4862]);
assign l_40[2799]    = ( l_41 [4863]);
assign l_40[2800]    = ( l_41 [4864]);
assign l_40[2801]    = ( l_41 [4865]);
assign l_40[2802]    = ( l_41 [4866]);
assign l_40[2803]    = ( l_41 [4867]);
assign l_40[2804]    = ( l_41 [4868]);
assign l_40[2805]    = ( l_41 [4869]);
assign l_40[2806]    = ( l_41 [4870]);
assign l_40[2807]    = ( l_41 [4871]);
assign l_40[2808]    = ( l_41 [4872]);
assign l_40[2809]    = ( l_41 [4873]);
assign l_40[2810]    = ( l_41 [4874]);
assign l_40[2811]    = ( l_41 [4875]);
assign l_40[2812]    = ( l_41 [4876]);
assign l_40[2813]    = ( l_41 [4877]);
assign l_40[2814]    = ( l_41 [4878]);
assign l_40[2815]    = ( l_41 [4879]);
assign l_40[2816]    = ( l_41 [4880]);
assign l_40[2817]    = ( l_41 [4881]);
assign l_40[2818]    = ( l_41 [4882]);
assign l_40[2819]    = ( l_41 [4883]);
assign l_40[2820]    = ( l_41 [4884]);
assign l_40[2821]    = ( l_41 [4885]);
assign l_40[2822]    = ( l_41 [4886]);
assign l_40[2823]    = ( l_41 [4887]);
assign l_40[2824]    = ( l_41 [4888]);
assign l_40[2825]    = ( l_41 [4889]);
assign l_40[2826]    = ( l_41 [4890]);
assign l_40[2827]    = ( l_41 [4891]);
assign l_40[2828]    = ( l_41 [4892]);
assign l_40[2829]    = ( l_41 [4893]);
assign l_40[2830]    = ( l_41 [4894]);
assign l_40[2831]    = ( l_41 [4895]);
assign l_40[2832]    = ( l_41 [4896]);
assign l_40[2833]    = ( l_41 [4897]);
assign l_40[2834]    = ( l_41 [4898]);
assign l_40[2835]    = ( l_41 [4899]);
assign l_40[2836]    = ( l_41 [4900]);
assign l_40[2837]    = ( l_41 [4901]);
assign l_40[2838]    = ( l_41 [4902]);
assign l_40[2839]    = ( l_41 [4903]);
assign l_40[2840]    = ( l_41 [4904]);
assign l_40[2841]    = ( l_41 [4905]);
assign l_40[2842]    = ( l_41 [4906]);
assign l_40[2843]    = ( l_41 [4907]);
assign l_40[2844]    = ( l_41 [4908]);
assign l_40[2845]    = ( l_41 [4909]);
assign l_40[2846]    = ( l_41 [4910]);
assign l_40[2847]    = ( l_41 [4911]);
assign l_40[2848]    = ( l_41 [4912]);
assign l_40[2849]    = ( l_41 [4913]);
assign l_40[2850]    = ( l_41 [4914]);
assign l_40[2851]    = ( l_41 [4915]);
assign l_40[2852]    = ( l_41 [4916]);
assign l_40[2853]    = ( l_41 [4917]);
assign l_40[2854]    = ( l_41 [4918]);
assign l_40[2855]    = ( l_41 [4919]);
assign l_40[2856]    = ( l_41 [4920]);
assign l_40[2857]    = ( l_41 [4921]);
assign l_40[2858]    = ( l_41 [4922]);
assign l_40[2859]    = ( l_41 [4923]);
assign l_40[2860]    = ( l_41 [4924]);
assign l_40[2861]    = ( l_41 [4925]);
assign l_40[2862]    = ( l_41 [4926]);
assign l_40[2863]    = ( l_41 [4927]);
assign l_40[2864]    = ( l_41 [4928]);
assign l_40[2865]    = ( l_41 [4929]);
assign l_40[2866]    = ( l_41 [4930]);
assign l_40[2867]    = ( l_41 [4931]);
assign l_40[2868]    = ( l_41 [4932]);
assign l_40[2869]    = ( l_41 [4933]);
assign l_40[2870]    = ( l_41 [4934]);
assign l_40[2871]    = ( l_41 [4935]);
assign l_40[2872]    = ( l_41 [4936]);
assign l_40[2873]    = ( l_41 [4937]);
assign l_40[2874]    = ( l_41 [4938]);
assign l_40[2875]    = ( l_41 [4939]);
assign l_40[2876]    = ( l_41 [4940]);
assign l_40[2877]    = ( l_41 [4941]);
assign l_40[2878]    = ( l_41 [4942]);
assign l_40[2879]    = ( l_41 [4943]);
assign l_40[2880]    = ( l_41 [4944]);
assign l_40[2881]    = ( l_41 [4945]);
assign l_40[2882]    = ( l_41 [4946]);
assign l_40[2883]    = ( l_41 [4947]);
assign l_40[2884]    = ( l_41 [4948]);
assign l_40[2885]    = ( l_41 [4949]);
assign l_40[2886]    = ( l_41 [4950]);
assign l_40[2887]    = ( l_41 [4951]);
assign l_40[2888]    = ( l_41 [4952]);
assign l_40[2889]    = ( l_41 [4953]);
assign l_40[2890]    = ( l_41 [4954]);
assign l_40[2891]    = ( l_41 [4955]);
assign l_40[2892]    = ( l_41 [4956]);
assign l_40[2893]    = ( l_41 [4957]);
assign l_40[2894]    = ( l_41 [4958]);
assign l_40[2895]    = ( l_41 [4959]);
assign l_40[2896]    = ( l_41 [4960]);
assign l_40[2897]    = ( l_41 [4961]);
assign l_40[2898]    = ( l_41 [4962]);
assign l_40[2899]    = ( l_41 [4963]);
assign l_40[2900]    = ( l_41 [4964]);
assign l_40[2901]    = ( l_41 [4965]);
assign l_40[2902]    = ( l_41 [4966]);
assign l_40[2903]    = ( l_41 [4967]);
assign l_40[2904]    = ( l_41 [4968]);
assign l_40[2905]    = ( l_41 [4969]);
assign l_40[2906]    = ( l_41 [4970]);
assign l_40[2907]    = ( l_41 [4971]);
assign l_40[2908]    = ( l_41 [4972]);
assign l_40[2909]    = ( l_41 [4973]);
assign l_40[2910]    = ( l_41 [4974]);
assign l_40[2911]    = ( l_41 [4975]);
assign l_40[2912]    = ( l_41 [4976]);
assign l_40[2913]    = ( l_41 [4977]);
assign l_40[2914]    = ( l_41 [4978]);
assign l_40[2915]    = ( l_41 [4979]);
assign l_40[2916]    = ( l_41 [4980]);
assign l_40[2917]    = ( l_41 [4981]);
assign l_40[2918]    = ( l_41 [4982]);
assign l_40[2919]    = ( l_41 [4983]);
assign l_40[2920]    = ( l_41 [4984]);
assign l_40[2921]    = ( l_41 [4985]);
assign l_40[2922]    = ( l_41 [4986]);
assign l_40[2923]    = ( l_41 [4987]);
assign l_40[2924]    = ( l_41 [4988]);
assign l_40[2925]    = ( l_41 [4989]);
assign l_40[2926]    = ( l_41 [4990]);
assign l_40[2927]    = ( l_41 [4991]);
assign l_40[2928]    = ( l_41 [4992]);
assign l_40[2929]    = ( l_41 [4993]);
assign l_40[2930]    = ( l_41 [4994]);
assign l_40[2931]    = ( l_41 [4995]);
assign l_40[2932]    = ( l_41 [4996]);
assign l_40[2933]    = ( l_41 [4997]);
assign l_40[2934]    = ( l_41 [4998]);
assign l_40[2935]    = ( l_41 [4999]);
assign l_40[2936]    = ( l_41 [5000]);
assign l_40[2937]    = ( l_41 [5001]);
assign l_40[2938]    = ( l_41 [5002]);
assign l_40[2939]    = ( l_41 [5003]);
assign l_40[2940]    = ( l_41 [5004]);
assign l_40[2941]    = ( l_41 [5005]);
assign l_40[2942]    = ( l_41 [5006]);
assign l_40[2943]    = ( l_41 [5007]);
assign l_40[2944]    = ( l_41 [5008]);
assign l_40[2945]    = ( l_41 [5009]);
assign l_40[2946]    = ( l_41 [5010]);
assign l_40[2947]    = ( l_41 [5011]);
assign l_40[2948]    = ( l_41 [5012]);
assign l_40[2949]    = ( l_41 [5013]);
assign l_40[2950]    = ( l_41 [5014]);
assign l_40[2951]    = ( l_41 [5015]);
assign l_40[2952]    = ( l_41 [5016]);
assign l_40[2953]    = ( l_41 [5017]);
assign l_40[2954]    = ( l_41 [5018]);
assign l_40[2955]    = ( l_41 [5019]);
assign l_40[2956]    = ( l_41 [5020]);
assign l_40[2957]    = ( l_41 [5021]);
assign l_40[2958]    = ( l_41 [5022]);
assign l_40[2959]    = ( l_41 [5023]);
assign l_40[2960]    = ( l_41 [5024]);
assign l_40[2961]    = ( l_41 [5025]);
assign l_40[2962]    = ( l_41 [5026]);
assign l_40[2963]    = ( l_41 [5027]);
assign l_40[2964]    = ( l_41 [5028]);
assign l_40[2965]    = ( l_41 [5029]);
assign l_40[2966]    = ( l_41 [5030]);
assign l_40[2967]    = ( l_41 [5031]);
assign l_40[2968]    = ( l_41 [5032]);
assign l_40[2969]    = ( l_41 [5033]);
assign l_40[2970]    = ( l_41 [5034]);
assign l_40[2971]    = ( l_41 [5035]);
assign l_40[2972]    = ( l_41 [5036]);
assign l_40[2973]    = ( l_41 [5037]);
assign l_40[2974]    = ( l_41 [5038]);
assign l_40[2975]    = ( l_41 [5039]);
assign l_40[2976]    = ( l_41 [5040]);
assign l_40[2977]    = ( l_41 [5041]);
assign l_40[2978]    = ( l_41 [5042]);
assign l_40[2979]    = ( l_41 [5043]);
assign l_40[2980]    = ( l_41 [5044]);
assign l_40[2981]    = ( l_41 [5045]);
assign l_40[2982]    = ( l_41 [5046]);
assign l_40[2983]    = ( l_41 [5047]);
assign l_40[2984]    = ( l_41 [5048]);
assign l_40[2985]    = ( l_41 [5049]);
assign l_40[2986]    = ( l_41 [5050]);
assign l_40[2987]    = ( l_41 [5051]);
assign l_40[2988]    = ( l_41 [5052]);
assign l_40[2989]    = ( l_41 [5053]);
assign l_40[2990]    = ( l_41 [5054]);
assign l_40[2991]    = ( l_41 [5055]);
assign l_40[2992]    = ( l_41 [5056]);
assign l_40[2993]    = ( l_41 [5057]);
assign l_40[2994]    = ( l_41 [5058]);
assign l_40[2995]    = ( l_41 [5059]);
assign l_40[2996]    = ( l_41 [5060]);
assign l_40[2997]    = ( l_41 [5061]);
assign l_40[2998]    = ( l_41 [5062]);
assign l_40[2999]    = ( l_41 [5063]);
assign l_40[3000]    = ( l_41 [5064]);
assign l_40[3001]    = ( l_41 [5065]);
assign l_40[3002]    = ( l_41 [5066]);
assign l_40[3003]    = ( l_41 [5067]);
assign l_40[3004]    = ( l_41 [5068]);
assign l_40[3005]    = ( l_41 [5069]);
assign l_40[3006]    = ( l_41 [5070]);
assign l_40[3007]    = ( l_41 [5071]);
assign l_40[3008]    = ( l_41 [5072]);
assign l_40[3009]    = ( l_41 [5073]);
assign l_40[3010]    = ( l_41 [5074]);
assign l_40[3011]    = ( l_41 [5075]);
assign l_40[3012]    = ( l_41 [5076]);
assign l_40[3013]    = ( l_41 [5077]);
assign l_40[3014]    = ( l_41 [5078]);
assign l_40[3015]    = ( l_41 [5079]);
assign l_40[3016]    = ( l_41 [5080]);
assign l_40[3017]    = ( l_41 [5081]);
assign l_40[3018]    = ( l_41 [5082]);
assign l_40[3019]    = ( l_41 [5083]);
assign l_40[3020]    = ( l_41 [5084]);
assign l_40[3021]    = ( l_41 [5085]);
assign l_40[3022]    = ( l_41 [5086]);
assign l_40[3023]    = ( l_41 [5087]);
assign l_40[3024]    = ( l_41 [5088]);
assign l_40[3025]    = ( l_41 [5089]);
assign l_40[3026]    = ( l_41 [5090]);
assign l_40[3027]    = ( l_41 [5091]);
assign l_40[3028]    = ( l_41 [5092]);
assign l_40[3029]    = ( l_41 [5093]);
assign l_40[3030]    = ( l_41 [5094]);
assign l_40[3031]    = ( l_41 [5095]);
assign l_40[3032]    = ( l_41 [5096]);
assign l_40[3033]    = ( l_41 [5097]);
assign l_40[3034]    = ( l_41 [5098]);
assign l_40[3035]    = ( l_41 [5099]);
assign l_40[3036]    = ( l_41 [5100]);
assign l_40[3037]    = ( l_41 [5101]);
assign l_40[3038]    = ( l_41 [5102]);
assign l_40[3039]    = ( l_41 [5103]);
assign l_40[3040]    = ( l_41 [5104]);
assign l_40[3041]    = ( l_41 [5105]);
assign l_40[3042]    = ( l_41 [5106]);
assign l_40[3043]    = ( l_41 [5107]);
assign l_40[3044]    = ( l_41 [5108]);
assign l_40[3045]    = ( l_41 [5109]);
assign l_40[3046]    = ( l_41 [5110]);
assign l_40[3047]    = ( l_41 [5111]);
assign l_40[3048]    = ( l_41 [5112]);
assign l_40[3049]    = ( l_41 [5113]);
assign l_40[3050]    = ( l_41 [5114]);
assign l_40[3051]    = ( l_41 [5115]);
assign l_40[3052]    = ( l_41 [5116]);
assign l_40[3053]    = ( l_41 [5117]);
assign l_40[3054]    = ( l_41 [5118]);
assign l_40[3055]    = ( l_41 [5119]);
assign l_40[3056]    = ( l_41 [5120]);
assign l_40[3057]    = ( l_41 [5121]);
assign l_40[3058]    = ( l_41 [5122]);
assign l_40[3059]    = ( l_41 [5123]);
assign l_40[3060]    = ( l_41 [5124]);
assign l_40[3061]    = ( l_41 [5125]);
assign l_40[3062]    = ( l_41 [5126]);
assign l_40[3063]    = ( l_41 [5127]);
assign l_40[3064]    = ( l_41 [5128]);
assign l_40[3065]    = ( l_41 [5129]);
assign l_40[3066]    = ( l_41 [5130]);
assign l_40[3067]    = ( l_41 [5131]);
assign l_40[3068]    = ( l_41 [5132]);
assign l_40[3069]    = ( l_41 [5133]);
assign l_40[3070]    = ( l_41 [5134]);
assign l_40[3071]    = ( l_41 [5135]);
assign l_40[3072]    = ( l_41 [5136]);
assign l_40[3073]    = ( l_41 [5137]);
assign l_40[3074]    = ( l_41 [5138]);
assign l_40[3075]    = ( l_41 [5139]);
assign l_40[3076]    = ( l_41 [5140]);
assign l_40[3077]    = ( l_41 [5141]);
assign l_40[3078]    = ( l_41 [5142]);
assign l_40[3079]    = ( l_41 [5143]);
assign l_40[3080]    = ( l_41 [5144]);
assign l_40[3081]    = ( l_41 [5145]);
assign l_40[3082]    = ( l_41 [5146]);
assign l_40[3083]    = ( l_41 [5147]);
assign l_40[3084]    = ( l_41 [5148]);
assign l_40[3085]    = ( l_41 [5149]);
assign l_40[3086]    = ( l_41 [5150]);
assign l_40[3087]    = ( l_41 [5151]);
assign l_40[3088]    = ( l_41 [5152]);
assign l_40[3089]    = ( l_41 [5153]);
assign l_40[3090]    = ( l_41 [5154]);
assign l_40[3091]    = ( l_41 [5155]);
assign l_40[3092]    = ( l_41 [5156]);
assign l_40[3093]    = ( l_41 [5157]);
assign l_40[3094]    = ( l_41 [5158]);
assign l_40[3095]    = ( l_41 [5159]);
assign l_40[3096]    = ( l_41 [5160]);
assign l_40[3097]    = ( l_41 [5161]);
assign l_40[3098]    = ( l_41 [5162]);
assign l_40[3099]    = ( l_41 [5163]);
assign l_40[3100]    = ( l_41 [5164]);
assign l_40[3101]    = ( l_41 [5165]);
assign l_40[3102]    = ( l_41 [5166]);
assign l_40[3103]    = ( l_41 [5167]);
assign l_40[3104]    = ( l_41 [5168]);
assign l_40[3105]    = ( l_41 [5169]);
assign l_40[3106]    = ( l_41 [5170]);
assign l_40[3107]    = ( l_41 [5171]);
assign l_40[3108]    = ( l_41 [5172]);
assign l_40[3109]    = ( l_41 [5173]);
assign l_40[3110]    = ( l_41 [5174]);
assign l_40[3111]    = ( l_41 [5175]);
assign l_40[3112]    = ( l_41 [5176]);
assign l_40[3113]    = ( l_41 [5177]);
assign l_40[3114]    = ( l_41 [5178]);
assign l_40[3115]    = ( l_41 [5179]);
assign l_40[3116]    = ( l_41 [5180]);
assign l_40[3117]    = ( l_41 [5181]);
assign l_40[3118]    = ( l_41 [5182]);
assign l_40[3119]    = ( l_41 [5183]);
assign l_40[3120]    = ( l_41 [5184]);
assign l_40[3121]    = ( l_41 [5185]);
assign l_40[3122]    = ( l_41 [5186]);
assign l_40[3123]    = ( l_41 [5187]);
assign l_40[3124]    = ( l_41 [5188]);
assign l_40[3125]    = ( l_41 [5189]);
assign l_40[3126]    = ( l_41 [5190]);
assign l_40[3127]    = ( l_41 [5191]);
assign l_40[3128]    = ( l_41 [5192]);
assign l_40[3129]    = ( l_41 [5193]);
assign l_40[3130]    = ( l_41 [5194]);
assign l_40[3131]    = ( l_41 [5195]);
assign l_40[3132]    = ( l_41 [5196]);
assign l_40[3133]    = ( l_41 [5197]);
assign l_40[3134]    = ( l_41 [5198]);
assign l_40[3135]    = ( l_41 [5199]);
assign l_40[3136]    = ( l_41 [5200]);
assign l_40[3137]    = ( l_41 [5201]);
assign l_40[3138]    = ( l_41 [5202]);
assign l_40[3139]    = ( l_41 [5203]);
assign l_40[3140]    = ( l_41 [5204]);
assign l_40[3141]    = ( l_41 [5205]);
assign l_40[3142]    = ( l_41 [5206]);
assign l_40[3143]    = ( l_41 [5207]);
assign l_40[3144]    = ( l_41 [5208]);
assign l_40[3145]    = ( l_41 [5209]);
assign l_40[3146]    = ( l_41 [5210]);
assign l_40[3147]    = ( l_41 [5211]);
assign l_40[3148]    = ( l_41 [5212]);
assign l_40[3149]    = ( l_41 [5213]);
assign l_40[3150]    = ( l_41 [5214]);
assign l_40[3151]    = ( l_41 [5215]);
assign l_40[3152]    = ( l_41 [5216]);
assign l_40[3153]    = ( l_41 [5217]);
assign l_40[3154]    = ( l_41 [5218]);
assign l_40[3155]    = ( l_41 [5219]);
assign l_40[3156]    = ( l_41 [5220]);
assign l_40[3157]    = ( l_41 [5221]);
assign l_40[3158]    = ( l_41 [5222]);
assign l_40[3159]    = ( l_41 [5223]);
assign l_40[3160]    = ( l_41 [5224]);
assign l_40[3161]    = ( l_41 [5225]);
assign l_40[3162]    = ( l_41 [5226]);
assign l_40[3163]    = ( l_41 [5227]);
assign l_40[3164]    = ( l_41 [5228]);
assign l_40[3165]    = ( l_41 [5229]);
assign l_40[3166]    = ( l_41 [5230]);
assign l_40[3167]    = ( l_41 [5231]);
assign l_40[3168]    = ( l_41 [5232]);
assign l_40[3169]    = ( l_41 [5233]);
assign l_40[3170]    = ( l_41 [5234]);
assign l_40[3171]    = ( l_41 [5235]);
assign l_40[3172]    = ( l_41 [5236]);
assign l_40[3173]    = ( l_41 [5237]);
assign l_40[3174]    = ( l_41 [5238]);
assign l_40[3175]    = ( l_41 [5239]);
assign l_40[3176]    = ( l_41 [5240]);
assign l_40[3177]    = ( l_41 [5241]);
assign l_40[3178]    = ( l_41 [5242]);
assign l_40[3179]    = ( l_41 [5243]);
assign l_40[3180]    = ( l_41 [5244]);
assign l_40[3181]    = ( l_41 [5245]);
assign l_40[3182]    = ( l_41 [5246]);
assign l_40[3183]    = ( l_41 [5247]);
assign l_40[3184]    = ( l_41 [5248]);
assign l_40[3185]    = ( l_41 [5249]);
assign l_40[3186]    = ( l_41 [5250]);
assign l_40[3187]    = ( l_41 [5251]);
assign l_40[3188]    = ( l_41 [5252]);
assign l_40[3189]    = ( l_41 [5253]);
assign l_40[3190]    = ( l_41 [5254]);
assign l_40[3191]    = ( l_41 [5255]);
assign l_40[3192]    = ( l_41 [5256]);
assign l_40[3193]    = ( l_41 [5257]);
assign l_40[3194]    = ( l_41 [5258]);
assign l_40[3195]    = ( l_41 [5259]);
assign l_40[3196]    = ( l_41 [5260]);
assign l_40[3197]    = ( l_41 [5261]);
assign l_40[3198]    = ( l_41 [5262]);
assign l_40[3199]    = ( l_41 [5263]);
assign l_40[3200]    = ( l_41 [5264]);
assign l_40[3201]    = ( l_41 [5265]);
assign l_40[3202]    = ( l_41 [5266]);
assign l_40[3203]    = ( l_41 [5267]);
assign l_40[3204]    = ( l_41 [5268]);
assign l_40[3205]    = ( l_41 [5269]);
assign l_40[3206]    = ( l_41 [5270]);
assign l_40[3207]    = ( l_41 [5271]);
assign l_40[3208]    = ( l_41 [5272]);
assign l_40[3209]    = ( l_41 [5273]);
assign l_40[3210]    = ( l_41 [5274]);
assign l_40[3211]    = ( l_41 [5275]);
assign l_40[3212]    = ( l_41 [5276]);
assign l_40[3213]    = ( l_41 [5277]);
assign l_40[3214]    = ( l_41 [5278]);
assign l_40[3215]    = ( l_41 [5279]);
assign l_40[3216]    = ( l_41 [5280]);
assign l_40[3217]    = ( l_41 [5281]);
assign l_40[3218]    = ( l_41 [5282]);
assign l_40[3219]    = ( l_41 [5283]);
assign l_40[3220]    = ( l_41 [5284]);
assign l_40[3221]    = ( l_41 [5285]);
assign l_40[3222]    = ( l_41 [5286]);
assign l_40[3223]    = ( l_41 [5287]);
assign l_40[3224]    = ( l_41 [5288]);
assign l_40[3225]    = ( l_41 [5289]);
assign l_40[3226]    = ( l_41 [5290]);
assign l_40[3227]    = ( l_41 [5291]);
assign l_40[3228]    = ( l_41 [5292]);
assign l_40[3229]    = ( l_41 [5293]);
assign l_40[3230]    = ( l_41 [5294]);
assign l_40[3231]    = ( l_41 [5295]);
assign l_40[3232]    = ( l_41 [5296]);
assign l_40[3233]    = ( l_41 [5297]);
assign l_40[3234]    = ( l_41 [5298]);
assign l_40[3235]    = ( l_41 [5299]);
assign l_40[3236]    = ( l_41 [5300]);
assign l_40[3237]    = ( l_41 [5301]);
assign l_40[3238]    = ( l_41 [5302]);
assign l_40[3239]    = ( l_41 [5303]);
assign l_40[3240]    = ( l_41 [5304]);
assign l_40[3241]    = ( l_41 [5305]);
assign l_40[3242]    = ( l_41 [5306]);
assign l_40[3243]    = ( l_41 [5307]);
assign l_40[3244]    = ( l_41 [5308]);
assign l_40[3245]    = ( l_41 [5309]);
assign l_40[3246]    = ( l_41 [5310]);
assign l_40[3247]    = ( l_41 [5311]);
assign l_40[3248]    = ( l_41 [5312]);
assign l_40[3249]    = ( l_41 [5313]);
assign l_40[3250]    = ( l_41 [5314]);
assign l_40[3251]    = ( l_41 [5315]);
assign l_40[3252]    = ( l_41 [5316]);
assign l_40[3253]    = ( l_41 [5317]);
assign l_40[3254]    = ( l_41 [5318]);
assign l_40[3255]    = ( l_41 [5319]);
assign l_40[3256]    = ( l_41 [5320]);
assign l_40[3257]    = ( l_41 [5321]);
assign l_40[3258]    = ( l_41 [5322]);
assign l_40[3259]    = ( l_41 [5323]);
assign l_40[3260]    = ( l_41 [5324]);
assign l_40[3261]    = ( l_41 [5325]);
assign l_40[3262]    = ( l_41 [5326]);
assign l_40[3263]    = ( l_41 [5327]);
assign l_40[3264]    = ( l_41 [5328]);
assign l_40[3265]    = ( l_41 [5329]);
assign l_40[3266]    = ( l_41 [5330]);
assign l_40[3267]    = ( l_41 [5331]);
assign l_40[3268]    = ( l_41 [5332]);
assign l_40[3269]    = ( l_41 [5333]);
assign l_40[3270]    = ( l_41 [5334]);
assign l_40[3271]    = ( l_41 [5335]);
assign l_40[3272]    = ( l_41 [5336]);
assign l_40[3273]    = ( l_41 [5337]);
assign l_40[3274]    = ( l_41 [5338]);
assign l_40[3275]    = ( l_41 [5339]);
assign l_40[3276]    = ( l_41 [5340]);
assign l_40[3277]    = ( l_41 [5341]);
assign l_40[3278]    = ( l_41 [5342]);
assign l_40[3279]    = ( l_41 [5343]);
assign l_40[3280]    = ( l_41 [5344]);
assign l_40[3281]    = ( l_41 [5345]);
assign l_40[3282]    = ( l_41 [5346]);
assign l_40[3283]    = ( l_41 [5347]);
assign l_40[3284]    = ( l_41 [5348]);
assign l_40[3285]    = ( l_41 [5349]);
assign l_40[3286]    = ( l_41 [5350]);
assign l_40[3287]    = ( l_41 [5351]);
assign l_40[3288]    = ( l_41 [5352]);
assign l_40[3289]    = ( l_41 [5353]);
assign l_40[3290]    = ( l_41 [5354]);
assign l_40[3291]    = ( l_41 [5355]);
assign l_40[3292]    = ( l_41 [5356]);
assign l_40[3293]    = ( l_41 [5357]);
assign l_40[3294]    = ( l_41 [5358]);
assign l_40[3295]    = ( l_41 [5359]);
assign l_40[3296]    = ( l_41 [5360]);
assign l_40[3297]    = ( l_41 [5361]);
assign l_40[3298]    = ( l_41 [5362]);
assign l_40[3299]    = ( l_41 [5363]);
assign l_40[3300]    = ( l_41 [5364]);
assign l_40[3301]    = ( l_41 [5365]);
assign l_40[3302]    = ( l_41 [5366]);
assign l_40[3303]    = ( l_41 [5367]);
assign l_40[3304]    = ( l_41 [5368]);
assign l_40[3305]    = ( l_41 [5369]);
assign l_40[3306]    = ( l_41 [5370]);
assign l_40[3307]    = ( l_41 [5371]);
assign l_40[3308]    = ( l_41 [5372]);
assign l_40[3309]    = ( l_41 [5373]);
assign l_40[3310]    = ( l_41 [5374]);
assign l_40[3311]    = ( l_41 [5375]);
assign l_40[3312]    = ( l_41 [5376]);
assign l_40[3313]    = ( l_41 [5377]);
assign l_40[3314]    = ( l_41 [5378]);
assign l_40[3315]    = ( l_41 [5379]);
assign l_40[3316]    = ( l_41 [5380]);
assign l_40[3317]    = ( l_41 [5381]);
assign l_40[3318]    = ( l_41 [5382]);
assign l_40[3319]    = ( l_41 [5383]);
assign l_40[3320]    = ( l_41 [5384]);
assign l_40[3321]    = ( l_41 [5385]);
assign l_40[3322]    = ( l_41 [5386]);
assign l_40[3323]    = ( l_41 [5387]);
assign l_40[3324]    = ( l_41 [5388]);
assign l_40[3325]    = ( l_41 [5389]);
assign l_40[3326]    = ( l_41 [5390]);
assign l_40[3327]    = ( l_41 [5391]);
assign l_40[3328]    = ( l_41 [5392]);
assign l_40[3329]    = ( l_41 [5393]);
assign l_40[3330]    = ( l_41 [5394]);
assign l_40[3331]    = ( l_41 [5395]);
assign l_40[3332]    = ( l_41 [5396]);
assign l_40[3333]    = ( l_41 [5397]);
assign l_40[3334]    = ( l_41 [5398]);
assign l_40[3335]    = ( l_41 [5399]);
assign l_40[3336]    = ( l_41 [5400]);
assign l_40[3337]    = ( l_41 [5401]);
assign l_40[3338]    = ( l_41 [5402]);
assign l_40[3339]    = ( l_41 [5403]);
assign l_40[3340]    = ( l_41 [5404]);
assign l_40[3341]    = ( l_41 [5405]);
assign l_40[3342]    = ( l_41 [5406]);
assign l_40[3343]    = ( l_41 [5407]);
assign l_40[3344]    = ( l_41 [5408]);
assign l_40[3345]    = ( l_41 [5409]);
assign l_40[3346]    = ( l_41 [5410]);
assign l_40[3347]    = ( l_41 [5411]);
assign l_40[3348]    = ( l_41 [5412]);
assign l_40[3349]    = ( l_41 [5413]);
assign l_40[3350]    = ( l_41 [5414]);
assign l_40[3351]    = ( l_41 [5415]);
assign l_40[3352]    = ( l_41 [5416]);
assign l_40[3353]    = ( l_41 [5417]);
assign l_40[3354]    = ( l_41 [5418]);
assign l_40[3355]    = ( l_41 [5419]);
assign l_40[3356]    = ( l_41 [5420]);
assign l_40[3357]    = ( l_41 [5421]);
assign l_40[3358]    = ( l_41 [5422]);
assign l_40[3359]    = ( l_41 [5423]);
assign l_40[3360]    = ( l_41 [5424]);
assign l_40[3361]    = ( l_41 [5425]);
assign l_40[3362]    = ( l_41 [5426]);
assign l_40[3363]    = ( l_41 [5427]);
assign l_40[3364]    = ( l_41 [5428]);
assign l_40[3365]    = ( l_41 [5429]);
assign l_40[3366]    = ( l_41 [5430]);
assign l_40[3367]    = ( l_41 [5431]);
assign l_40[3368]    = ( l_41 [5432]);
assign l_40[3369]    = ( l_41 [5433]);
assign l_40[3370]    = ( l_41 [5434]);
assign l_40[3371]    = ( l_41 [5435]);
assign l_40[3372]    = ( l_41 [5436]);
assign l_40[3373]    = ( l_41 [5437]);
assign l_40[3374]    = ( l_41 [5438]);
assign l_40[3375]    = ( l_41 [5439]);
assign l_40[3376]    = ( l_41 [5440]);
assign l_40[3377]    = ( l_41 [5441]);
assign l_40[3378]    = ( l_41 [5442]);
assign l_40[3379]    = ( l_41 [5443]);
assign l_40[3380]    = ( l_41 [5444]);
assign l_40[3381]    = ( l_41 [5445]);
assign l_40[3382]    = ( l_41 [5446]);
assign l_40[3383]    = ( l_41 [5447]);
assign l_40[3384]    = ( l_41 [5448]);
assign l_40[3385]    = ( l_41 [5449]);
assign l_40[3386]    = ( l_41 [5450]);
assign l_40[3387]    = ( l_41 [5451]);
assign l_40[3388]    = ( l_41 [5452]);
assign l_40[3389]    = ( l_41 [5453]);
assign l_40[3390]    = ( l_41 [5454]);
assign l_40[3391]    = ( l_41 [5455]);
assign l_40[3392]    = ( l_41 [5456]);
assign l_40[3393]    = ( l_41 [5457]);
assign l_40[3394]    = ( l_41 [5458]);
assign l_40[3395]    = ( l_41 [5459]);
assign l_40[3396]    = ( l_41 [5460]);
assign l_40[3397]    = ( l_41 [5461]);
assign l_40[3398]    = ( l_41 [5462]);
assign l_40[3399]    = ( l_41 [5463]);
assign l_40[3400]    = ( l_41 [5464]);
assign l_40[3401]    = ( l_41 [5465]);
assign l_40[3402]    = ( l_41 [5466]);
assign l_40[3403]    = ( l_41 [5467]);
assign l_40[3404]    = ( l_41 [5468]);
assign l_40[3405]    = ( l_41 [5469]);
assign l_40[3406]    = ( l_41 [5470]);
assign l_40[3407]    = ( l_41 [5471]);
assign l_40[3408]    = ( l_41 [5472]);
assign l_40[3409]    = ( l_41 [5473]);
assign l_40[3410]    = ( l_41 [5474]);
assign l_40[3411]    = ( l_41 [5475]);
assign l_40[3412]    = ( l_41 [5476]);
assign l_40[3413]    = ( l_41 [5477]);
assign l_40[3414]    = ( l_41 [5478]);
assign l_40[3415]    = ( l_41 [5479]);
assign l_40[3416]    = ( l_41 [5480]);
assign l_40[3417]    = ( l_41 [5481]);
assign l_40[3418]    = ( l_41 [5482]);
assign l_40[3419]    = ( l_41 [5483]);
assign l_40[3420]    = ( l_41 [5484]);
assign l_40[3421]    = ( l_41 [5485]);
assign l_40[3422]    = ( l_41 [5486]);
assign l_40[3423]    = ( l_41 [5487]);
assign l_40[3424]    = ( l_41 [5488]);
assign l_40[3425]    = ( l_41 [5489]);
assign l_40[3426]    = ( l_41 [5490]);
assign l_40[3427]    = ( l_41 [5491]);
assign l_40[3428]    = ( l_41 [5492]);
assign l_40[3429]    = ( l_41 [5493]);
assign l_40[3430]    = ( l_41 [5494]);
assign l_40[3431]    = ( l_41 [5495]);
assign l_40[3432]    = ( l_41 [5496]);
assign l_40[3433]    = ( l_41 [5497]);
assign l_40[3434]    = ( l_41 [5498]);
assign l_40[3435]    = ( l_41 [5499]);
assign l_40[3436]    = ( l_41 [5500]);
assign l_40[3437]    = ( l_41 [5501]);
assign l_40[3438]    = ( l_41 [5502]);
assign l_40[3439]    = ( l_41 [5503]);
assign l_40[3440]    = ( l_41 [5504]);
assign l_40[3441]    = ( l_41 [5505]);
assign l_40[3442]    = ( l_41 [5506]);
assign l_40[3443]    = ( l_41 [5507]);
assign l_40[3444]    = ( l_41 [5508]);
assign l_40[3445]    = ( l_41 [5509]);
assign l_40[3446]    = ( l_41 [5510]);
assign l_40[3447]    = ( l_41 [5511]);
assign l_40[3448]    = ( l_41 [5512]);
assign l_40[3449]    = ( l_41 [5513]);
assign l_40[3450]    = ( l_41 [5514]);
assign l_40[3451]    = ( l_41 [5515]);
assign l_40[3452]    = ( l_41 [5516]);
assign l_40[3453]    = ( l_41 [5517]);
assign l_40[3454]    = ( l_41 [5518]);
assign l_40[3455]    = ( l_41 [5519]);
assign l_40[3456]    = ( l_41 [5520]);
assign l_40[3457]    = ( l_41 [5521]);
assign l_40[3458]    = ( l_41 [5522]);
assign l_40[3459]    = ( l_41 [5523]);
assign l_40[3460]    = ( l_41 [5524]);
assign l_40[3461]    = ( l_41 [5525]);
assign l_40[3462]    = ( l_41 [5526]);
assign l_40[3463]    = ( l_41 [5527]);
assign l_40[3464]    = ( l_41 [5528]);
assign l_40[3465]    = ( l_41 [5529]);
assign l_40[3466]    = ( l_41 [5530]);
assign l_40[3467]    = ( l_41 [5531]);
assign l_40[3468]    = ( l_41 [5532]);
assign l_40[3469]    = ( l_41 [5533]);
assign l_40[3470]    = ( l_41 [5534]);
assign l_40[3471]    = ( l_41 [5535]);
assign l_40[3472]    = ( l_41 [5536]);
assign l_40[3473]    = ( l_41 [5537]);
assign l_40[3474]    = ( l_41 [5538]);
assign l_40[3475]    = ( l_41 [5539]);
assign l_40[3476]    = ( l_41 [5540]);
assign l_40[3477]    = ( l_41 [5541]);
assign l_40[3478]    = ( l_41 [5542]);
assign l_40[3479]    = ( l_41 [5543]);
assign l_40[3480]    = ( l_41 [5544]);
assign l_40[3481]    = ( l_41 [5545]);
assign l_40[3482]    = ( l_41 [5546]);
assign l_40[3483]    = ( l_41 [5547]);
assign l_40[3484]    = ( l_41 [5548]);
assign l_40[3485]    = ( l_41 [5549]);
assign l_40[3486]    = ( l_41 [5550]);
assign l_40[3487]    = ( l_41 [5551]);
assign l_40[3488]    = ( l_41 [5552]);
assign l_40[3489]    = ( l_41 [5553]);
assign l_40[3490]    = ( l_41 [5554]);
assign l_40[3491]    = ( l_41 [5555]);
assign l_40[3492]    = ( l_41 [5556]);
assign l_40[3493]    = ( l_41 [5557]);
assign l_40[3494]    = ( l_41 [5558]);
assign l_40[3495]    = ( l_41 [5559]);
assign l_40[3496]    = ( l_41 [5560]);
assign l_40[3497]    = ( l_41 [5561]);
assign l_40[3498]    = ( l_41 [5562]);
assign l_40[3499]    = ( l_41 [5563]);
assign l_40[3500]    = ( l_41 [5564]);
assign l_40[3501]    = ( l_41 [5565]);
assign l_40[3502]    = ( l_41 [5566]);
assign l_40[3503]    = ( l_41 [5567]);
assign l_40[3504]    = ( l_41 [5568]);
assign l_40[3505]    = ( l_41 [5569]);
assign l_40[3506]    = ( l_41 [5570]);
assign l_40[3507]    = ( l_41 [5571]);
assign l_40[3508]    = ( l_41 [5572]);
assign l_40[3509]    = ( l_41 [5573]);
assign l_40[3510]    = ( l_41 [5574]);
assign l_40[3511]    = ( l_41 [5575]);
assign l_40[3512]    = ( l_41 [5576]);
assign l_40[3513]    = ( l_41 [5577]);
assign l_40[3514]    = ( l_41 [5578]);
assign l_40[3515]    = ( l_41 [5579]);
assign l_40[3516]    = ( l_41 [5580]);
assign l_40[3517]    = ( l_41 [5581]);
assign l_40[3518]    = ( l_41 [5582]);
assign l_40[3519]    = ( l_41 [5583]);
assign l_40[3520]    = ( l_41 [5584]);
assign l_40[3521]    = ( l_41 [5585]);
assign l_40[3522]    = ( l_41 [5586]);
assign l_40[3523]    = ( l_41 [5587]);
assign l_40[3524]    = ( l_41 [5588]);
assign l_40[3525]    = ( l_41 [5589]);
assign l_40[3526]    = ( l_41 [5590]);
assign l_40[3527]    = ( l_41 [5591]);
assign l_40[3528]    = ( l_41 [5592]);
assign l_40[3529]    = ( l_41 [5593]);
assign l_40[3530]    = ( l_41 [5594]);
assign l_40[3531]    = ( l_41 [5595]);
assign l_40[3532]    = ( l_41 [5596]);
assign l_40[3533]    = ( l_41 [5597]);
assign l_40[3534]    = ( l_41 [5598]);
assign l_40[3535]    = ( l_41 [5599]);
assign l_40[3536]    = ( l_41 [5600]);
assign l_40[3537]    = ( l_41 [5601]);
assign l_40[3538]    = ( l_41 [5602]);
assign l_40[3539]    = ( l_41 [5603]);
assign l_40[3540]    = ( l_41 [5604]);
assign l_40[3541]    = ( l_41 [5605]);
assign l_40[3542]    = ( l_41 [5606]);
assign l_40[3543]    = ( l_41 [5607]);
assign l_40[3544]    = ( l_41 [5608]);
assign l_40[3545]    = ( l_41 [5609]);
assign l_40[3546]    = ( l_41 [5610]);
assign l_40[3547]    = ( l_41 [5611]);
assign l_40[3548]    = ( l_41 [5612]);
assign l_40[3549]    = ( l_41 [5613]);
assign l_40[3550]    = ( l_41 [5614]);
assign l_40[3551]    = ( l_41 [5615]);
assign l_40[3552]    = ( l_41 [5616]);
assign l_40[3553]    = ( l_41 [5617]);
assign l_40[3554]    = ( l_41 [5618]);
assign l_40[3555]    = ( l_41 [5619]);
assign l_40[3556]    = ( l_41 [5620]);
assign l_40[3557]    = ( l_41 [5621]);
assign l_40[3558]    = ( l_41 [5622]);
assign l_40[3559]    = ( l_41 [5623]);
assign l_40[3560]    = ( l_41 [5624]);
assign l_40[3561]    = ( l_41 [5625]);
assign l_40[3562]    = ( l_41 [5626]);
assign l_40[3563]    = ( l_41 [5627]);
assign l_40[3564]    = ( l_41 [5628]);
assign l_40[3565]    = ( l_41 [5629]);
assign l_40[3566]    = ( l_41 [5630]);
assign l_40[3567]    = ( l_41 [5631]);
assign l_40[3568]    = ( l_41 [5632]);
assign l_40[3569]    = ( l_41 [5633]);
assign l_40[3570]    = ( l_41 [5634]);
assign l_40[3571]    = ( l_41 [5635]);
assign l_40[3572]    = ( l_41 [5636]);
assign l_40[3573]    = ( l_41 [5637]);
assign l_40[3574]    = ( l_41 [5638]);
assign l_40[3575]    = ( l_41 [5639]);
assign l_40[3576]    = ( l_41 [5640]);
assign l_40[3577]    = ( l_41 [5641]);
assign l_40[3578]    = ( l_41 [5642]);
assign l_40[3579]    = ( l_41 [5643]);
assign l_40[3580]    = ( l_41 [5644]);
assign l_40[3581]    = ( l_41 [5645]);
assign l_40[3582]    = ( l_41 [5646]);
assign l_40[3583]    = ( l_41 [5647]);
assign l_40[3584]    = ( l_41 [5648]);
assign l_40[3585]    = ( l_41 [5649]);
assign l_40[3586]    = ( l_41 [5650]);
assign l_40[3587]    = ( l_41 [5651]);
assign l_40[3588]    = ( l_41 [5652]);
assign l_40[3589]    = ( l_41 [5653]);
assign l_40[3590]    = ( l_41 [5654]);
assign l_40[3591]    = ( l_41 [5655]);
assign l_40[3592]    = ( l_41 [5656]);
assign l_40[3593]    = ( l_41 [5657]);
assign l_40[3594]    = ( l_41 [5658]);
assign l_40[3595]    = ( l_41 [5659]);
assign l_40[3596]    = ( l_41 [5660]);
assign l_40[3597]    = ( l_41 [5661]);
assign l_40[3598]    = ( l_41 [5662]);
assign l_40[3599]    = ( l_41 [5663]);
assign l_40[3600]    = ( l_41 [5664]);
assign l_40[3601]    = ( l_41 [5665]);
assign l_40[3602]    = ( l_41 [5666]);
assign l_40[3603]    = ( l_41 [5667]);
assign l_40[3604]    = ( l_41 [5668]);
assign l_40[3605]    = ( l_41 [5669]);
assign l_40[3606]    = ( l_41 [5670]);
assign l_40[3607]    = ( l_41 [5671]);
assign l_40[3608]    = ( l_41 [5672]);
assign l_40[3609]    = ( l_41 [5673]);
assign l_40[3610]    = ( l_41 [5674]);
assign l_40[3611]    = ( l_41 [5675]);
assign l_40[3612]    = ( l_41 [5676]);
assign l_40[3613]    = ( l_41 [5677]);
assign l_40[3614]    = ( l_41 [5678]);
assign l_40[3615]    = ( l_41 [5679]);
assign l_40[3616]    = ( l_41 [5680]);
assign l_40[3617]    = ( l_41 [5681]);
assign l_40[3618]    = ( l_41 [5682]);
assign l_40[3619]    = ( l_41 [5683]);
assign l_40[3620]    = ( l_41 [5684]);
assign l_40[3621]    = ( l_41 [5685]);
assign l_40[3622]    = ( l_41 [5686]);
assign l_40[3623]    = ( l_41 [5687]);
assign l_40[3624]    = ( l_41 [5688]);
assign l_40[3625]    = ( l_41 [5689]);
assign l_40[3626]    = ( l_41 [5690]);
assign l_40[3627]    = ( l_41 [5691]);
assign l_40[3628]    = ( l_41 [5692]);
assign l_40[3629]    = ( l_41 [5693]);
assign l_40[3630]    = ( l_41 [5694]);
assign l_40[3631]    = ( l_41 [5695]);
assign l_40[3632]    = ( l_41 [5696]);
assign l_40[3633]    = ( l_41 [5697]);
assign l_40[3634]    = ( l_41 [5698]);
assign l_40[3635]    = ( l_41 [5699]);
assign l_40[3636]    = ( l_41 [5700]);
assign l_40[3637]    = ( l_41 [5701]);
assign l_40[3638]    = ( l_41 [5702]);
assign l_40[3639]    = ( l_41 [5703]);
assign l_40[3640]    = ( l_41 [5704]);
assign l_40[3641]    = ( l_41 [5705]);
assign l_40[3642]    = ( l_41 [5706]);
assign l_40[3643]    = ( l_41 [5707]);
assign l_40[3644]    = ( l_41 [5708]);
assign l_40[3645]    = ( l_41 [5709]);
assign l_40[3646]    = ( l_41 [5710]);
assign l_40[3647]    = ( l_41 [5711]);
assign l_40[3648]    = ( l_41 [5712]);
assign l_40[3649]    = ( l_41 [5713]);
assign l_40[3650]    = ( l_41 [5714]);
assign l_40[3651]    = ( l_41 [5715]);
assign l_40[3652]    = ( l_41 [5716]);
assign l_40[3653]    = ( l_41 [5717]);
assign l_40[3654]    = ( l_41 [5718]);
assign l_40[3655]    = ( l_41 [5719]);
assign l_40[3656]    = ( l_41 [5720]);
assign l_40[3657]    = ( l_41 [5721]);
assign l_40[3658]    = ( l_41 [5722]);
assign l_40[3659]    = ( l_41 [5723]);
assign l_40[3660]    = ( l_41 [5724]);
assign l_40[3661]    = ( l_41 [5725]);
assign l_40[3662]    = ( l_41 [5726]);
assign l_40[3663]    = ( l_41 [5727]);
assign l_40[3664]    = ( l_41 [5728]);
assign l_40[3665]    = ( l_41 [5729]);
assign l_40[3666]    = ( l_41 [5730]);
assign l_40[3667]    = ( l_41 [5731]);
assign l_40[3668]    = ( l_41 [5732]);
assign l_40[3669]    = ( l_41 [5733]);
assign l_40[3670]    = ( l_41 [5734]);
assign l_40[3671]    = ( l_41 [5735]);
assign l_40[3672]    = ( l_41 [5736]);
assign l_40[3673]    = ( l_41 [5737]);
assign l_40[3674]    = ( l_41 [5738]);
assign l_40[3675]    = ( l_41 [5739]);
assign l_40[3676]    = ( l_41 [5740]);
assign l_40[3677]    = ( l_41 [5741]);
assign l_40[3678]    = ( l_41 [5742]);
assign l_40[3679]    = ( l_41 [5743]);
assign l_40[3680]    = ( l_41 [5744]);
assign l_40[3681]    = ( l_41 [5745]);
assign l_40[3682]    = ( l_41 [5746]);
assign l_40[3683]    = ( l_41 [5747]);
assign l_40[3684]    = ( l_41 [5748]);
assign l_40[3685]    = ( l_41 [5749]);
assign l_40[3686]    = ( l_41 [5750]);
assign l_40[3687]    = ( l_41 [5751]);
assign l_40[3688]    = ( l_41 [5752]);
assign l_40[3689]    = ( l_41 [5753]);
assign l_40[3690]    = ( l_41 [5754]);
assign l_40[3691]    = ( l_41 [5755]);
assign l_40[3692]    = ( l_41 [5756]);
assign l_40[3693]    = ( l_41 [5757]);
assign l_40[3694]    = ( l_41 [5758]);
assign l_40[3695]    = ( l_41 [5759]);
assign l_40[3696]    = ( l_41 [5760]);
assign l_40[3697]    = ( l_41 [5761]);
assign l_40[3698]    = ( l_41 [5762]);
assign l_40[3699]    = ( l_41 [5763]);
assign l_40[3700]    = ( l_41 [5764]);
assign l_40[3701]    = ( l_41 [5765]);
assign l_40[3702]    = ( l_41 [5766]);
assign l_40[3703]    = ( l_41 [5767]);
assign l_40[3704]    = ( l_41 [5768]);
assign l_40[3705]    = ( l_41 [5769]);
assign l_40[3706]    = ( l_41 [5770]);
assign l_40[3707]    = ( l_41 [5771]);
assign l_40[3708]    = ( l_41 [5772]);
assign l_40[3709]    = ( l_41 [5773]);
assign l_40[3710]    = ( l_41 [5774]);
assign l_40[3711]    = ( l_41 [5775]);
assign l_40[3712]    = ( l_41 [5776]);
assign l_40[3713]    = ( l_41 [5777]);
assign l_40[3714]    = ( l_41 [5778]);
assign l_40[3715]    = ( l_41 [5779]);
assign l_40[3716]    = ( l_41 [5780]);
assign l_40[3717]    = ( l_41 [5781]);
assign l_40[3718]    = ( l_41 [5782]);
assign l_40[3719]    = ( l_41 [5783]);
assign l_40[3720]    = ( l_41 [5784]);
assign l_40[3721]    = ( l_41 [5785]);
assign l_40[3722]    = ( l_41 [5786]);
assign l_40[3723]    = ( l_41 [5787]);
assign l_40[3724]    = ( l_41 [5788]);
assign l_40[3725]    = ( l_41 [5789]);
assign l_40[3726]    = ( l_41 [5790]);
assign l_40[3727]    = ( l_41 [5791]);
assign l_40[3728]    = ( l_41 [5792]);
assign l_40[3729]    = ( l_41 [5793]);
assign l_40[3730]    = ( l_41 [5794]);
assign l_40[3731]    = ( l_41 [5795]);
assign l_40[3732]    = ( l_41 [5796]);
assign l_40[3733]    = ( l_41 [5797]);
assign l_40[3734]    = ( l_41 [5798]);
assign l_40[3735]    = ( l_41 [5799]);
assign l_40[3736]    = ( l_41 [5800]);
assign l_40[3737]    = ( l_41 [5801]);
assign l_40[3738]    = ( l_41 [5802]);
assign l_40[3739]    = ( l_41 [5803]);
assign l_40[3740]    = ( l_41 [5804]);
assign l_40[3741]    = ( l_41 [5805]);
assign l_40[3742]    = ( l_41 [5806]);
assign l_40[3743]    = ( l_41 [5807]);
assign l_40[3744]    = ( l_41 [5808]);
assign l_40[3745]    = ( l_41 [5809]);
assign l_40[3746]    = ( l_41 [5810]);
assign l_40[3747]    = ( l_41 [5811]);
assign l_40[3748]    = ( l_41 [5812]);
assign l_40[3749]    = ( l_41 [5813]);
assign l_40[3750]    = ( l_41 [5814]);
assign l_40[3751]    = ( l_41 [5815]);
assign l_40[3752]    = ( l_41 [5816]);
assign l_40[3753]    = ( l_41 [5817]);
assign l_40[3754]    = ( l_41 [5818]);
assign l_40[3755]    = ( l_41 [5819]);
assign l_40[3756]    = ( l_41 [5820]);
assign l_40[3757]    = ( l_41 [5821]);
assign l_40[3758]    = ( l_41 [5822]);
assign l_40[3759]    = ( l_41 [5823]);
assign l_40[3760]    = ( l_41 [5824]);
assign l_40[3761]    = ( l_41 [5825]);
assign l_40[3762]    = ( l_41 [5826]);
assign l_40[3763]    = ( l_41 [5827]);
assign l_40[3764]    = ( l_41 [5828]);
assign l_40[3765]    = ( l_41 [5829]);
assign l_40[3766]    = ( l_41 [5830]);
assign l_40[3767]    = ( l_41 [5831]);
assign l_40[3768]    = ( l_41 [5832]);
assign l_40[3769]    = ( l_41 [5833]);
assign l_40[3770]    = ( l_41 [5834]);
assign l_40[3771]    = ( l_41 [5835]);
assign l_40[3772]    = ( l_41 [5836]);
assign l_40[3773]    = ( l_41 [5837]);
assign l_40[3774]    = ( l_41 [5838]);
assign l_40[3775]    = ( l_41 [5839]);
assign l_40[3776]    = ( l_41 [5840]);
assign l_40[3777]    = ( l_41 [5841]);
assign l_40[3778]    = ( l_41 [5842]);
assign l_40[3779]    = ( l_41 [5843]);
assign l_40[3780]    = ( l_41 [5844]);
assign l_40[3781]    = ( l_41 [5845]);
assign l_40[3782]    = ( l_41 [5846]);
assign l_40[3783]    = ( l_41 [5847]);
assign l_40[3784]    = ( l_41 [5848]);
assign l_40[3785]    = ( l_41 [5849]);
assign l_40[3786]    = ( l_41 [5850]);
assign l_40[3787]    = ( l_41 [5851]);
assign l_40[3788]    = ( l_41 [5852]);
assign l_40[3789]    = ( l_41 [5853]);
assign l_40[3790]    = ( l_41 [5854]);
assign l_40[3791]    = ( l_41 [5855]);
assign l_40[3792]    = ( l_41 [5856]);
assign l_40[3793]    = ( l_41 [5857]);
assign l_40[3794]    = ( l_41 [5858]);
assign l_40[3795]    = ( l_41 [5859]);
assign l_40[3796]    = ( l_41 [5860]);
assign l_40[3797]    = ( l_41 [5861]);
assign l_40[3798]    = ( l_41 [5862]);
assign l_40[3799]    = ( l_41 [5863]);
assign l_40[3800]    = ( l_41 [5864]);
assign l_40[3801]    = ( l_41 [5865]);
assign l_40[3802]    = ( l_41 [5866]);
assign l_40[3803]    = ( l_41 [5867]);
assign l_40[3804]    = ( l_41 [5868]);
assign l_40[3805]    = ( l_41 [5869]);
assign l_40[3806]    = ( l_41 [5870]);
assign l_40[3807]    = ( l_41 [5871]);
assign l_40[3808]    = ( l_41 [5872]);
assign l_40[3809]    = ( l_41 [5873]);
assign l_40[3810]    = ( l_41 [5874]);
assign l_40[3811]    = ( l_41 [5875]);
assign l_40[3812]    = ( l_41 [5876]);
assign l_40[3813]    = ( l_41 [5877]);
assign l_40[3814]    = ( l_41 [5878]);
assign l_40[3815]    = ( l_41 [5879]);
assign l_40[3816]    = ( l_41 [5880]);
assign l_40[3817]    = ( l_41 [5881]);
assign l_40[3818]    = ( l_41 [5882]);
assign l_40[3819]    = ( l_41 [5883]);
assign l_40[3820]    = ( l_41 [5884]);
assign l_40[3821]    = ( l_41 [5885]);
assign l_40[3822]    = ( l_41 [5886]);
assign l_40[3823]    = ( l_41 [5887]);
assign l_40[3824]    = ( l_41 [5888]);
assign l_40[3825]    = ( l_41 [5889]);
assign l_40[3826]    = ( l_41 [5890]);
assign l_40[3827]    = ( l_41 [5891]);
assign l_40[3828]    = ( l_41 [5892]);
assign l_40[3829]    = ( l_41 [5893]);
assign l_40[3830]    = ( l_41 [5894]);
assign l_40[3831]    = ( l_41 [5895]);
assign l_40[3832]    = ( l_41 [5896]);
assign l_40[3833]    = ( l_41 [5897]);
assign l_40[3834]    = ( l_41 [5898]);
assign l_40[3835]    = ( l_41 [5899]);
assign l_40[3836]    = ( l_41 [5900]);
assign l_40[3837]    = ( l_41 [5901]);
assign l_40[3838]    = ( l_41 [5902]);
assign l_40[3839]    = ( l_41 [5903]);
assign l_40[3840]    = ( l_41 [5904]);
assign l_40[3841]    = ( l_41 [5905]);
assign l_40[3842]    = ( l_41 [5906]);
assign l_40[3843]    = ( l_41 [5907]);
assign l_40[3844]    = ( l_41 [5908]);
assign l_40[3845]    = ( l_41 [5909]);
assign l_40[3846]    = ( l_41 [5910]);
assign l_40[3847]    = ( l_41 [5911]);
assign l_40[3848]    = ( l_41 [5912]);
assign l_40[3849]    = ( l_41 [5913]);
assign l_40[3850]    = ( l_41 [5914]);
assign l_40[3851]    = ( l_41 [5915]);
assign l_40[3852]    = ( l_41 [5916]);
assign l_40[3853]    = ( l_41 [5917]);
assign l_40[3854]    = ( l_41 [5918]);
assign l_40[3855]    = ( l_41 [5919]);
assign l_40[3856]    = ( l_41 [5920]);
assign l_40[3857]    = ( l_41 [5921]);
assign l_40[3858]    = ( l_41 [5922]);
assign l_40[3859]    = ( l_41 [5923]);
assign l_40[3860]    = ( l_41 [5924]);
assign l_40[3861]    = ( l_41 [5925]);
assign l_40[3862]    = ( l_41 [5926]);
assign l_40[3863]    = ( l_41 [5927]);
assign l_40[3864]    = ( l_41 [5928]);
assign l_40[3865]    = ( l_41 [5929]);
assign l_40[3866]    = ( l_41 [5930]);
assign l_40[3867]    = ( l_41 [5931]);
assign l_40[3868]    = ( l_41 [5932]);
assign l_40[3869]    = ( l_41 [5933]);
assign l_40[3870]    = ( l_41 [5934]);
assign l_40[3871]    = ( l_41 [5935]);
assign l_40[3872]    = ( l_41 [5936]);
assign l_40[3873]    = ( l_41 [5937]);
assign l_40[3874]    = ( l_41 [5938]);
assign l_40[3875]    = ( l_41 [5939]);
assign l_40[3876]    = ( l_41 [5940]);
assign l_40[3877]    = ( l_41 [5941]);
assign l_40[3878]    = ( l_41 [5942]);
assign l_40[3879]    = ( l_41 [5943]);
assign l_40[3880]    = ( l_41 [5944]);
assign l_40[3881]    = ( l_41 [5945]);
assign l_40[3882]    = ( l_41 [5946]);
assign l_40[3883]    = ( l_41 [5947]);
assign l_40[3884]    = ( l_41 [5948]);
assign l_40[3885]    = ( l_41 [5949]);
assign l_40[3886]    = ( l_41 [5950]);
assign l_40[3887]    = ( l_41 [5951]);
assign l_40[3888]    = ( l_41 [5952]);
assign l_40[3889]    = ( l_41 [5953]);
assign l_40[3890]    = ( l_41 [5954]);
assign l_40[3891]    = ( l_41 [5955]);
assign l_40[3892]    = ( l_41 [5956]);
assign l_40[3893]    = ( l_41 [5957]);
assign l_40[3894]    = ( l_41 [5958]);
assign l_40[3895]    = ( l_41 [5959]);
assign l_40[3896]    = ( l_41 [5960]);
assign l_40[3897]    = ( l_41 [5961]);
assign l_40[3898]    = ( l_41 [5962]);
assign l_40[3899]    = ( l_41 [5963]);
assign l_40[3900]    = ( l_41 [5964]);
assign l_40[3901]    = ( l_41 [5965]);
assign l_40[3902]    = ( l_41 [5966]);
assign l_40[3903]    = ( l_41 [5967]);
assign l_40[3904]    = ( l_41 [5968]);
assign l_40[3905]    = ( l_41 [5969]);
assign l_40[3906]    = ( l_41 [5970]);
assign l_40[3907]    = ( l_41 [5971]);
assign l_40[3908]    = ( l_41 [5972]);
assign l_40[3909]    = ( l_41 [5973]);
assign l_40[3910]    = ( l_41 [5974]);
assign l_40[3911]    = ( l_41 [5975]);
assign l_40[3912]    = ( l_41 [5976]);
assign l_40[3913]    = ( l_41 [5977]);
assign l_40[3914]    = ( l_41 [5978]);
assign l_40[3915]    = ( l_41 [5979]);
assign l_40[3916]    = ( l_41 [5980]);
assign l_40[3917]    = ( l_41 [5981]);
assign l_40[3918]    = ( l_41 [5982]);
assign l_40[3919]    = ( l_41 [5983]);
assign l_40[3920]    = ( l_41 [5984]);
assign l_40[3921]    = ( l_41 [5985]);
assign l_40[3922]    = ( l_41 [5986]);
assign l_40[3923]    = ( l_41 [5987]);
assign l_40[3924]    = ( l_41 [5988]);
assign l_40[3925]    = ( l_41 [5989]);
assign l_40[3926]    = ( l_41 [5990]);
assign l_40[3927]    = ( l_41 [5991]);
assign l_40[3928]    = ( l_41 [5992]);
assign l_40[3929]    = ( l_41 [5993]);
assign l_40[3930]    = ( l_41 [5994]);
assign l_40[3931]    = ( l_41 [5995]);
assign l_40[3932]    = ( l_41 [5996]);
assign l_40[3933]    = ( l_41 [5997]);
assign l_40[3934]    = ( l_41 [5998]);
assign l_40[3935]    = ( l_41 [5999]);
assign l_40[3936]    = ( l_41 [6000]);
assign l_40[3937]    = ( l_41 [6001]);
assign l_40[3938]    = ( l_41 [6002]);
assign l_40[3939]    = ( l_41 [6003]);
assign l_40[3940]    = ( l_41 [6004]);
assign l_40[3941]    = ( l_41 [6005]);
assign l_40[3942]    = ( l_41 [6006]);
assign l_40[3943]    = ( l_41 [6007]);
assign l_40[3944]    = ( l_41 [6008]);
assign l_40[3945]    = ( l_41 [6009]);
assign l_40[3946]    = ( l_41 [6010]);
assign l_40[3947]    = ( l_41 [6011]);
assign l_40[3948]    = ( l_41 [6012]);
assign l_40[3949]    = ( l_41 [6013]);
assign l_40[3950]    = ( l_41 [6014]);
assign l_40[3951]    = ( l_41 [6015]);
assign l_40[3952]    = ( l_41 [6016]);
assign l_40[3953]    = ( l_41 [6017]);
assign l_40[3954]    = ( l_41 [6018]);
assign l_40[3955]    = ( l_41 [6019]);
assign l_40[3956]    = ( l_41 [6020]);
assign l_40[3957]    = ( l_41 [6021]);
assign l_40[3958]    = ( l_41 [6022]);
assign l_40[3959]    = ( l_41 [6023]);
assign l_40[3960]    = ( l_41 [6024]);
assign l_40[3961]    = ( l_41 [6025]);
assign l_40[3962]    = ( l_41 [6026]);
assign l_40[3963]    = ( l_41 [6027]);
assign l_40[3964]    = ( l_41 [6028]);
assign l_40[3965]    = ( l_41 [6029]);
assign l_40[3966]    = ( l_41 [6030]);
assign l_40[3967]    = ( l_41 [6031]);
assign l_40[3968]    = ( l_41 [6032]);
assign l_40[3969]    = ( l_41 [6033]);
assign l_40[3970]    = ( l_41 [6034]);
assign l_40[3971]    = ( l_41 [6035]);
assign l_40[3972]    = ( l_41 [6036]);
assign l_40[3973]    = ( l_41 [6037]);
assign l_40[3974]    = ( l_41 [6038]);
assign l_40[3975]    = ( l_41 [6039]);
assign l_40[3976]    = ( l_41 [6040]);
assign l_40[3977]    = ( l_41 [6041]);
assign l_40[3978]    = ( l_41 [6042]);
assign l_40[3979]    = ( l_41 [6043]);
assign l_40[3980]    = ( l_41 [6044]);
assign l_40[3981]    = ( l_41 [6045]);
assign l_40[3982]    = ( l_41 [6046]);
assign l_40[3983]    = ( l_41 [6047]);
assign l_40[3984]    = ( l_41 [6048]);
assign l_40[3985]    = ( l_41 [6049]);
assign l_40[3986]    = ( l_41 [6050]);
assign l_40[3987]    = ( l_41 [6051]);
assign l_40[3988]    = ( l_41 [6052]);
assign l_40[3989]    = ( l_41 [6053]);
assign l_40[3990]    = ( l_41 [6054]);
assign l_40[3991]    = ( l_41 [6055]);
assign l_40[3992]    = ( l_41 [6056]);
assign l_40[3993]    = ( l_41 [6057]);
assign l_40[3994]    = ( l_41 [6058]);
assign l_40[3995]    = ( l_41 [6059]);
assign l_40[3996]    = ( l_41 [6060]);
assign l_40[3997]    = ( l_41 [6061]);
assign l_40[3998]    = ( l_41 [6062]);
assign l_40[3999]    = ( l_41 [6063]);
assign l_40[4000]    = ( l_41 [6064]);
assign l_40[4001]    = ( l_41 [6065]);
assign l_40[4002]    = ( l_41 [6066]);
assign l_40[4003]    = ( l_41 [6067]);
assign l_40[4004]    = ( l_41 [6068]);
assign l_40[4005]    = ( l_41 [6069]);
assign l_40[4006]    = ( l_41 [6070]);
assign l_40[4007]    = ( l_41 [6071]);
assign l_40[4008]    = ( l_41 [6072]);
assign l_40[4009]    = ( l_41 [6073]);
assign l_40[4010]    = ( l_41 [6074]);
assign l_40[4011]    = ( l_41 [6075]);
assign l_40[4012]    = ( l_41 [6076]);
assign l_40[4013]    = ( l_41 [6077]);
assign l_40[4014]    = ( l_41 [6078]);
assign l_40[4015]    = ( l_41 [6079]);
assign l_40[4016]    = ( l_41 [6080]);
assign l_40[4017]    = ( l_41 [6081]);
assign l_40[4018]    = ( l_41 [6082]);
assign l_40[4019]    = ( l_41 [6083]);
assign l_40[4020]    = ( l_41 [6084]);
assign l_40[4021]    = ( l_41 [6085]);
assign l_40[4022]    = ( l_41 [6086]);
assign l_40[4023]    = ( l_41 [6087]);
assign l_40[4024]    = ( l_41 [6088]);
assign l_40[4025]    = ( l_41 [6089]);
assign l_40[4026]    = ( l_41 [6090]);
assign l_40[4027]    = ( l_41 [6091]);
assign l_40[4028]    = ( l_41 [6092]);
assign l_40[4029]    = ( l_41 [6093]);
assign l_40[4030]    = ( l_41 [6094]);
assign l_40[4031]    = ( l_41 [6095]);
assign l_40[4032]    = ( l_41 [6096]);
assign l_40[4033]    = ( l_41 [6097]);
assign l_40[4034]    = ( l_41 [6098]);
assign l_40[4035]    = ( l_41 [6099]);
assign l_40[4036]    = ( l_41 [6100]);
assign l_40[4037]    = ( l_41 [6101]);
assign l_40[4038]    = ( l_41 [6102]);
assign l_40[4039]    = ( l_41 [6103]);
assign l_40[4040]    = ( l_41 [6104]);
assign l_40[4041]    = ( l_41 [6105]);
assign l_40[4042]    = ( l_41 [6106]);
assign l_40[4043]    = ( l_41 [6107]);
assign l_40[4044]    = ( l_41 [6108]);
assign l_40[4045]    = ( l_41 [6109]);
assign l_40[4046]    = ( l_41 [6110]);
assign l_40[4047]    = ( l_41 [6111]);
assign l_40[4048]    = ( l_41 [6112]);
assign l_40[4049]    = ( l_41 [6113]);
assign l_40[4050]    = ( l_41 [6114]);
assign l_40[4051]    = ( l_41 [6115]);
assign l_40[4052]    = ( l_41 [6116]);
assign l_40[4053]    = ( l_41 [6117]);
assign l_40[4054]    = ( l_41 [6118]);
assign l_40[4055]    = ( l_41 [6119]);
assign l_40[4056]    = ( l_41 [6120]);
assign l_40[4057]    = ( l_41 [6121]);
assign l_40[4058]    = ( l_41 [6122]);
assign l_40[4059]    = ( l_41 [6123]);
assign l_40[4060]    = ( l_41 [6124]);
assign l_40[4061]    = ( l_41 [6125]);
assign l_40[4062]    = ( l_41 [6126]);
assign l_40[4063]    = ( l_41 [6127]);
assign l_40[4064]    = ( l_41 [6128]);
assign l_40[4065]    = ( l_41 [6129]);
assign l_40[4066]    = ( l_41 [6130]);
assign l_40[4067]    = ( l_41 [6131]);
assign l_40[4068]    = ( l_41 [6132]);
assign l_40[4069]    = ( l_41 [6133]);
assign l_40[4070]    = ( l_41 [6134]);
assign l_40[4071]    = ( l_41 [6135]);
assign l_40[4072]    = ( l_41 [6136]);
assign l_40[4073]    = ( l_41 [6137]);
assign l_40[4074]    = ( l_41 [6138]);
assign l_40[4075]    = ( l_41 [6139]);
assign l_40[4076]    = ( l_41 [6140]);
assign l_40[4077]    = ( l_41 [6141]);
assign l_40[4078]    = ( l_41 [6142]);
assign l_40[4079]    = ( l_41 [6143]);
assign l_40[4080]    = ( l_41 [6144]);
assign l_40[4081]    = ( l_41 [6145]);
assign l_40[4082]    = ( l_41 [6146]);
assign l_40[4083]    = ( l_41 [6147]);
assign l_40[4084]    = ( l_41 [6148]);
assign l_40[4085]    = ( l_41 [6149]);
assign l_40[4086]    = ( l_41 [6150]);
assign l_40[4087]    = ( l_41 [6151]);
assign l_40[4088]    = ( l_41 [6152]);
assign l_40[4089]    = ( l_41 [6153]);
assign l_40[4090]    = ( l_41 [6154]);
assign l_40[4091]    = ( l_41 [6155]);
assign l_40[4092]    = ( l_41 [6156]);
assign l_40[4093]    = ( l_41 [6157]);
assign l_40[4094]    = ( l_41 [6158]);
assign l_40[4095]    = ( l_41 [6159]);
assign l_40[4096]    = ( l_41 [6160]);
assign l_40[4097]    = ( l_41 [6161]);
assign l_40[4098]    = ( l_41 [6162]);
assign l_40[4099]    = ( l_41 [6163]);
assign l_40[4100]    = ( l_41 [6164]);
assign l_40[4101]    = ( l_41 [6165]);
assign l_40[4102]    = ( l_41 [6166]);
assign l_40[4103]    = ( l_41 [6167]);
assign l_40[4104]    = ( l_41 [6168]);
assign l_40[4105]    = ( l_41 [6169]);
assign l_40[4106]    = ( l_41 [6170]);
assign l_40[4107]    = ( l_41 [6171]);
assign l_40[4108]    = ( l_41 [6172]);
assign l_40[4109]    = ( l_41 [6173]);
assign l_40[4110]    = ( l_41 [6174]);
assign l_40[4111]    = ( l_41 [6175]);
assign l_40[4112]    = ( l_41 [6176]);
assign l_40[4113]    = ( l_41 [6177]);
assign l_41[0]    = ( l_42 [0]);
assign l_41[1]    = ( l_42 [1] & !i[1820]) | ( l_42 [2] &  i[1820]);
assign l_41[2]    = ( l_42 [3] & !i[1820]) | ( l_42 [4] &  i[1820]);
assign l_41[3]    = ( l_42 [5] & !i[1820]) | ( l_42 [6] &  i[1820]);
assign l_41[4]    = ( l_42 [7] & !i[1820]) | ( l_42 [8] &  i[1820]);
assign l_41[5]    = ( l_42 [9] & !i[1820]) | ( l_42 [10] &  i[1820]);
assign l_41[6]    = ( l_42 [11] & !i[1820]) | ( l_42 [12] &  i[1820]);
assign l_41[7]    = ( l_42 [13] & !i[1820]) | ( l_42 [14] &  i[1820]);
assign l_41[8]    = ( l_42 [15] & !i[1820]) | ( l_42 [16] &  i[1820]);
assign l_41[9]    = ( l_42 [17] & !i[1820]) | ( l_42 [18] &  i[1820]);
assign l_41[10]    = ( l_42 [19] & !i[1820]) | ( l_42 [20] &  i[1820]);
assign l_41[11]    = ( l_42 [21] & !i[1820]) | ( l_42 [22] &  i[1820]);
assign l_41[12]    = ( l_42 [23] & !i[1820]) | ( l_42 [24] &  i[1820]);
assign l_41[13]    = ( l_42 [25] & !i[1820]) | ( l_42 [26] &  i[1820]);
assign l_41[14]    = ( l_42 [27] & !i[1820]) | ( l_42 [28] &  i[1820]);
assign l_41[15]    = ( l_42 [29] & !i[1820]) | ( l_42 [30] &  i[1820]);
assign l_41[16]    = ( l_42 [31] & !i[1820]) | ( l_42 [32] &  i[1820]);
assign l_41[17]    = ( l_42 [33] & !i[1820]) | ( l_42 [34] &  i[1820]);
assign l_41[18]    = ( l_42 [35] & !i[1820]) | ( l_42 [36] &  i[1820]);
assign l_41[19]    = ( l_42 [37]);
assign l_41[20]    = ( l_42 [38] & !i[1820]) | ( l_42 [39] &  i[1820]);
assign l_41[21]    = ( l_42 [40] & !i[1820]) | ( l_42 [41] &  i[1820]);
assign l_41[22]    = ( l_42 [42] & !i[1820]) | ( l_42 [43] &  i[1820]);
assign l_41[23]    = ( l_42 [44] & !i[1820]) | ( l_42 [45] &  i[1820]);
assign l_41[24]    = ( l_42 [46] & !i[1820]) | ( l_42 [47] &  i[1820]);
assign l_41[25]    = ( l_42 [48] & !i[1820]) | ( l_42 [49] &  i[1820]);
assign l_41[26]    = ( l_42 [50] & !i[1820]) | ( l_42 [51] &  i[1820]);
assign l_41[27]    = ( l_42 [52] & !i[1820]) | ( l_42 [53] &  i[1820]);
assign l_41[28]    = ( l_42 [54] & !i[1820]) | ( l_42 [55] &  i[1820]);
assign l_41[29]    = ( l_42 [56] & !i[1820]) | ( l_42 [57] &  i[1820]);
assign l_41[30]    = ( l_42 [58] & !i[1820]) | ( l_42 [59] &  i[1820]);
assign l_41[31]    = ( l_42 [60] & !i[1820]) | ( l_42 [61] &  i[1820]);
assign l_41[32]    = ( l_42 [62] & !i[1820]) | ( l_42 [63] &  i[1820]);
assign l_41[33]    = ( l_42 [64] & !i[1820]) | ( l_42 [65] &  i[1820]);
assign l_41[34]    = ( l_42 [66]);
assign l_41[35]    = ( l_42 [67]);
assign l_41[36]    = ( l_42 [68]);
assign l_41[37]    = ( l_42 [69]);
assign l_41[38]    = ( l_42 [70]);
assign l_41[39]    = ( l_42 [71]);
assign l_41[40]    = ( l_42 [72]);
assign l_41[41]    = ( l_42 [73]);
assign l_41[42]    = ( l_42 [74]);
assign l_41[43]    = ( l_42 [75]);
assign l_41[44]    = ( l_42 [76]);
assign l_41[45]    = ( l_42 [77]);
assign l_41[46]    = ( l_42 [78]);
assign l_41[47]    = ( l_42 [79]);
assign l_41[48]    = ( l_42 [80]);
assign l_41[49]    = ( l_42 [81]);
assign l_41[50]    = ( l_42 [82]);
assign l_41[51]    = ( l_42 [83]);
assign l_41[52]    = ( l_42 [84]);
assign l_41[53]    = ( l_42 [85]);
assign l_41[54]    = ( l_42 [86]);
assign l_41[55]    = ( l_42 [87]);
assign l_41[56]    = ( l_42 [88]);
assign l_41[57]    = ( l_42 [89]);
assign l_41[58]    = ( l_42 [90]);
assign l_41[59]    = ( l_42 [91]);
assign l_41[60]    = ( l_42 [92]);
assign l_41[61]    = ( l_42 [93]);
assign l_41[62]    = ( l_42 [94]);
assign l_41[63]    = ( l_42 [95]);
assign l_41[64]    = ( l_42 [96]);
assign l_41[65]    = ( l_42 [97]);
assign l_41[66]    = ( l_42 [98]);
assign l_41[67]    = ( l_42 [99]);
assign l_41[68]    = ( l_42 [100]);
assign l_41[69]    = ( l_42 [101]);
assign l_41[70]    = ( l_42 [102]);
assign l_41[71]    = ( l_42 [103]);
assign l_41[72]    = ( l_42 [104]);
assign l_41[73]    = ( l_42 [105]);
assign l_41[74]    = ( l_42 [106]);
assign l_41[75]    = ( l_42 [107]);
assign l_41[76]    = ( l_42 [108]);
assign l_41[77]    = ( l_42 [109]);
assign l_41[78]    = ( l_42 [110]);
assign l_41[79]    = ( l_42 [111]);
assign l_41[80]    = ( l_42 [112]);
assign l_41[81]    = ( l_42 [113]);
assign l_41[82]    = ( l_42 [114]);
assign l_41[83]    = ( l_42 [115]);
assign l_41[84]    = ( l_42 [116]);
assign l_41[85]    = ( l_42 [117]);
assign l_41[86]    = ( l_42 [118]);
assign l_41[87]    = ( l_42 [119]);
assign l_41[88]    = ( l_42 [120]);
assign l_41[89]    = ( l_42 [121]);
assign l_41[90]    = ( l_42 [122]);
assign l_41[91]    = ( l_42 [123]);
assign l_41[92]    = ( l_42 [124]);
assign l_41[93]    = ( l_42 [125]);
assign l_41[94]    = ( l_42 [126]);
assign l_41[95]    = ( l_42 [127]);
assign l_41[96]    = ( l_42 [128]);
assign l_41[97]    = ( l_42 [129]);
assign l_41[98]    = ( l_42 [130]);
assign l_41[99]    = ( l_42 [131]);
assign l_41[100]    = ( l_42 [132]);
assign l_41[101]    = ( l_42 [133]);
assign l_41[102]    = ( l_42 [134]);
assign l_41[103]    = ( l_42 [135]);
assign l_41[104]    = ( l_42 [136]);
assign l_41[105]    = ( l_42 [137]);
assign l_41[106]    = ( l_42 [138]);
assign l_41[107]    = ( l_42 [139]);
assign l_41[108]    = ( l_42 [140]);
assign l_41[109]    = ( l_42 [141]);
assign l_41[110]    = ( l_42 [142]);
assign l_41[111]    = ( l_42 [143]);
assign l_41[112]    = ( l_42 [144]);
assign l_41[113]    = ( l_42 [145]);
assign l_41[114]    = ( l_42 [146]);
assign l_41[115]    = ( l_42 [147]);
assign l_41[116]    = ( l_42 [148]);
assign l_41[117]    = ( l_42 [149]);
assign l_41[118]    = ( l_42 [150]);
assign l_41[119]    = ( l_42 [151]);
assign l_41[120]    = ( l_42 [152]);
assign l_41[121]    = ( l_42 [153]);
assign l_41[122]    = ( l_42 [154]);
assign l_41[123]    = ( l_42 [155]);
assign l_41[124]    = ( l_42 [156]);
assign l_41[125]    = ( l_42 [157]);
assign l_41[126]    = ( l_42 [158]);
assign l_41[127]    = ( l_42 [159]);
assign l_41[128]    = ( l_42 [160]);
assign l_41[129]    = ( l_42 [161]);
assign l_41[130]    = ( l_42 [162]);
assign l_41[131]    = ( l_42 [163]);
assign l_41[132]    = ( l_42 [164]);
assign l_41[133]    = ( l_42 [165]);
assign l_41[134]    = ( l_42 [166]);
assign l_41[135]    = ( l_42 [167]);
assign l_41[136]    = ( l_42 [168]);
assign l_41[137]    = ( l_42 [169]);
assign l_41[138]    = ( l_42 [170]);
assign l_41[139]    = ( l_42 [171]);
assign l_41[140]    = ( l_42 [172]);
assign l_41[141]    = ( l_42 [173]);
assign l_41[142]    = ( l_42 [174]);
assign l_41[143]    = ( l_42 [175]);
assign l_41[144]    = ( l_42 [176]);
assign l_41[145]    = ( l_42 [177]);
assign l_41[146]    = ( l_42 [178]);
assign l_41[147]    = ( l_42 [179]);
assign l_41[148]    = ( l_42 [180]);
assign l_41[149]    = ( l_42 [181]);
assign l_41[150]    = ( l_42 [182]);
assign l_41[151]    = ( l_42 [183]);
assign l_41[152]    = ( l_42 [184]);
assign l_41[153]    = ( l_42 [185]);
assign l_41[154]    = ( l_42 [186]);
assign l_41[155]    = ( l_42 [187]);
assign l_41[156]    = ( l_42 [188]);
assign l_41[157]    = ( l_42 [189]);
assign l_41[158]    = ( l_42 [190]);
assign l_41[159]    = ( l_42 [191]);
assign l_41[160]    = ( l_42 [192]);
assign l_41[161]    = ( l_42 [193]);
assign l_41[162]    = ( l_42 [194]);
assign l_41[163]    = ( l_42 [195]);
assign l_41[164]    = ( l_42 [196]);
assign l_41[165]    = ( l_42 [197]);
assign l_41[166]    = ( l_42 [198]);
assign l_41[167]    = ( l_42 [199]);
assign l_41[168]    = ( l_42 [200]);
assign l_41[169]    = ( l_42 [201]);
assign l_41[170]    = ( l_42 [202]);
assign l_41[171]    = ( l_42 [203]);
assign l_41[172]    = ( l_42 [204]);
assign l_41[173]    = ( l_42 [205]);
assign l_41[174]    = ( l_42 [206]);
assign l_41[175]    = ( l_42 [207]);
assign l_41[176]    = ( l_42 [208]);
assign l_41[177]    = ( l_42 [209]);
assign l_41[178]    = ( l_42 [210]);
assign l_41[179]    = ( l_42 [211]);
assign l_41[180]    = ( l_42 [212]);
assign l_41[181]    = ( l_42 [213]);
assign l_41[182]    = ( l_42 [214]);
assign l_41[183]    = ( l_42 [215]);
assign l_41[184]    = ( l_42 [216]);
assign l_41[185]    = ( l_42 [217]);
assign l_41[186]    = ( l_42 [218]);
assign l_41[187]    = ( l_42 [219]);
assign l_41[188]    = ( l_42 [220]);
assign l_41[189]    = ( l_42 [221]);
assign l_41[190]    = ( l_42 [222]);
assign l_41[191]    = ( l_42 [223]);
assign l_41[192]    = ( l_42 [224]);
assign l_41[193]    = ( l_42 [225]);
assign l_41[194]    = ( l_42 [226]);
assign l_41[195]    = ( l_42 [227]);
assign l_41[196]    = ( l_42 [228]);
assign l_41[197]    = ( l_42 [229]);
assign l_41[198]    = ( l_42 [230]);
assign l_41[199]    = ( l_42 [231]);
assign l_41[200]    = ( l_42 [232]);
assign l_41[201]    = ( l_42 [233]);
assign l_41[202]    = ( l_42 [234]);
assign l_41[203]    = ( l_42 [235]);
assign l_41[204]    = ( l_42 [236]);
assign l_41[205]    = ( l_42 [237]);
assign l_41[206]    = ( l_42 [238]);
assign l_41[207]    = ( l_42 [239]);
assign l_41[208]    = ( l_42 [240]);
assign l_41[209]    = ( l_42 [241]);
assign l_41[210]    = ( l_42 [242]);
assign l_41[211]    = ( l_42 [243]);
assign l_41[212]    = ( l_42 [244]);
assign l_41[213]    = ( l_42 [245]);
assign l_41[214]    = ( l_42 [246]);
assign l_41[215]    = ( l_42 [247]);
assign l_41[216]    = ( l_42 [248]);
assign l_41[217]    = ( l_42 [249]);
assign l_41[218]    = ( l_42 [250]);
assign l_41[219]    = ( l_42 [251]);
assign l_41[220]    = ( l_42 [252]);
assign l_41[221]    = ( l_42 [253]);
assign l_41[222]    = ( l_42 [254]);
assign l_41[223]    = ( l_42 [255]);
assign l_41[224]    = ( l_42 [256]);
assign l_41[225]    = ( l_42 [257]);
assign l_41[226]    = ( l_42 [258]);
assign l_41[227]    = ( l_42 [259]);
assign l_41[228]    = ( l_42 [260]);
assign l_41[229]    = ( l_42 [261]);
assign l_41[230]    = ( l_42 [262]);
assign l_41[231]    = ( l_42 [263]);
assign l_41[232]    = ( l_42 [264]);
assign l_41[233]    = ( l_42 [265]);
assign l_41[234]    = ( l_42 [266]);
assign l_41[235]    = ( l_42 [267]);
assign l_41[236]    = ( l_42 [268]);
assign l_41[237]    = ( l_42 [269]);
assign l_41[238]    = ( l_42 [270]);
assign l_41[239]    = ( l_42 [271]);
assign l_41[240]    = ( l_42 [272]);
assign l_41[241]    = ( l_42 [273]);
assign l_41[242]    = ( l_42 [274]);
assign l_41[243]    = ( l_42 [275]);
assign l_41[244]    = ( l_42 [276]);
assign l_41[245]    = ( l_42 [277]);
assign l_41[246]    = ( l_42 [278]);
assign l_41[247]    = ( l_42 [279]);
assign l_41[248]    = ( l_42 [280]);
assign l_41[249]    = ( l_42 [281]);
assign l_41[250]    = ( l_42 [282]);
assign l_41[251]    = ( l_42 [283]);
assign l_41[252]    = ( l_42 [284]);
assign l_41[253]    = ( l_42 [285]);
assign l_41[254]    = ( l_42 [286]);
assign l_41[255]    = ( l_42 [287]);
assign l_41[256]    = ( l_42 [288]);
assign l_41[257]    = ( l_42 [289]);
assign l_41[258]    = ( l_42 [290]);
assign l_41[259]    = ( l_42 [291]);
assign l_41[260]    = ( l_42 [292]);
assign l_41[261]    = ( l_42 [293]);
assign l_41[262]    = ( l_42 [294]);
assign l_41[263]    = ( l_42 [295]);
assign l_41[264]    = ( l_42 [296]);
assign l_41[265]    = ( l_42 [297]);
assign l_41[266]    = ( l_42 [298]);
assign l_41[267]    = ( l_42 [299]);
assign l_41[268]    = ( l_42 [300]);
assign l_41[269]    = ( l_42 [301]);
assign l_41[270]    = ( l_42 [302]);
assign l_41[271]    = ( l_42 [303]);
assign l_41[272]    = ( l_42 [304]);
assign l_41[273]    = ( l_42 [305]);
assign l_41[274]    = ( l_42 [306]);
assign l_41[275]    = ( l_42 [307]);
assign l_41[276]    = ( l_42 [308]);
assign l_41[277]    = ( l_42 [309]);
assign l_41[278]    = ( l_42 [310]);
assign l_41[279]    = ( l_42 [311]);
assign l_41[280]    = ( l_42 [312]);
assign l_41[281]    = ( l_42 [313]);
assign l_41[282]    = ( l_42 [314]);
assign l_41[283]    = ( l_42 [315]);
assign l_41[284]    = ( l_42 [316]);
assign l_41[285]    = ( l_42 [317]);
assign l_41[286]    = ( l_42 [318]);
assign l_41[287]    = ( l_42 [319]);
assign l_41[288]    = ( l_42 [320]);
assign l_41[289]    = ( l_42 [321]);
assign l_41[290]    = ( l_42 [322]);
assign l_41[291]    = ( l_42 [323]);
assign l_41[292]    = ( l_42 [324]);
assign l_41[293]    = ( l_42 [325]);
assign l_41[294]    = ( l_42 [326]);
assign l_41[295]    = ( l_42 [327]);
assign l_41[296]    = ( l_42 [328]);
assign l_41[297]    = ( l_42 [329]);
assign l_41[298]    = ( l_42 [330]);
assign l_41[299]    = ( l_42 [331]);
assign l_41[300]    = ( l_42 [332]);
assign l_41[301]    = ( l_42 [333]);
assign l_41[302]    = ( l_42 [334]);
assign l_41[303]    = ( l_42 [335]);
assign l_41[304]    = ( l_42 [336]);
assign l_41[305]    = ( l_42 [337]);
assign l_41[306]    = ( l_42 [338]);
assign l_41[307]    = ( l_42 [339]);
assign l_41[308]    = ( l_42 [340]);
assign l_41[309]    = ( l_42 [341]);
assign l_41[310]    = ( l_42 [342]);
assign l_41[311]    = ( l_42 [343]);
assign l_41[312]    = ( l_42 [344]);
assign l_41[313]    = ( l_42 [345]);
assign l_41[314]    = ( l_42 [346]);
assign l_41[315]    = ( l_42 [347]);
assign l_41[316]    = ( l_42 [348]);
assign l_41[317]    = ( l_42 [349]);
assign l_41[318]    = ( l_42 [350]);
assign l_41[319]    = ( l_42 [351]);
assign l_41[320]    = ( l_42 [352]);
assign l_41[321]    = ( l_42 [353]);
assign l_41[322]    = ( l_42 [354]);
assign l_41[323]    = ( l_42 [355]);
assign l_41[324]    = ( l_42 [356]);
assign l_41[325]    = ( l_42 [357]);
assign l_41[326]    = ( l_42 [358]);
assign l_41[327]    = ( l_42 [359]);
assign l_41[328]    = ( l_42 [360]);
assign l_41[329]    = ( l_42 [361]);
assign l_41[330]    = ( l_42 [362]);
assign l_41[331]    = ( l_42 [363]);
assign l_41[332]    = ( l_42 [364]);
assign l_41[333]    = ( l_42 [365]);
assign l_41[334]    = ( l_42 [366]);
assign l_41[335]    = ( l_42 [367]);
assign l_41[336]    = ( l_42 [368]);
assign l_41[337]    = ( l_42 [369]);
assign l_41[338]    = ( l_42 [370]);
assign l_41[339]    = ( l_42 [371]);
assign l_41[340]    = ( l_42 [372]);
assign l_41[341]    = ( l_42 [373]);
assign l_41[342]    = ( l_42 [374]);
assign l_41[343]    = ( l_42 [375]);
assign l_41[344]    = ( l_42 [376]);
assign l_41[345]    = ( l_42 [377]);
assign l_41[346]    = ( l_42 [378]);
assign l_41[347]    = ( l_42 [379]);
assign l_41[348]    = ( l_42 [380]);
assign l_41[349]    = ( l_42 [381]);
assign l_41[350]    = ( l_42 [382]);
assign l_41[351]    = ( l_42 [383]);
assign l_41[352]    = ( l_42 [384]);
assign l_41[353]    = ( l_42 [385]);
assign l_41[354]    = ( l_42 [386]);
assign l_41[355]    = ( l_42 [387]);
assign l_41[356]    = ( l_42 [388]);
assign l_41[357]    = ( l_42 [389]);
assign l_41[358]    = ( l_42 [390]);
assign l_41[359]    = ( l_42 [391]);
assign l_41[360]    = ( l_42 [392]);
assign l_41[361]    = ( l_42 [393]);
assign l_41[362]    = ( l_42 [394]);
assign l_41[363]    = ( l_42 [395]);
assign l_41[364]    = ( l_42 [396]);
assign l_41[365]    = ( l_42 [397]);
assign l_41[366]    = ( l_42 [398]);
assign l_41[367]    = ( l_42 [399]);
assign l_41[368]    = ( l_42 [400]);
assign l_41[369]    = ( l_42 [401]);
assign l_41[370]    = ( l_42 [402]);
assign l_41[371]    = ( l_42 [403]);
assign l_41[372]    = ( l_42 [404]);
assign l_41[373]    = ( l_42 [405]);
assign l_41[374]    = ( l_42 [406]);
assign l_41[375]    = ( l_42 [407]);
assign l_41[376]    = ( l_42 [408]);
assign l_41[377]    = ( l_42 [409]);
assign l_41[378]    = ( l_42 [410]);
assign l_41[379]    = ( l_42 [411]);
assign l_41[380]    = ( l_42 [412]);
assign l_41[381]    = ( l_42 [413]);
assign l_41[382]    = ( l_42 [414]);
assign l_41[383]    = ( l_42 [415]);
assign l_41[384]    = ( l_42 [416]);
assign l_41[385]    = ( l_42 [417]);
assign l_41[386]    = ( l_42 [418]);
assign l_41[387]    = ( l_42 [419]);
assign l_41[388]    = ( l_42 [420]);
assign l_41[389]    = ( l_42 [421]);
assign l_41[390]    = ( l_42 [422]);
assign l_41[391]    = ( l_42 [423]);
assign l_41[392]    = ( l_42 [424]);
assign l_41[393]    = ( l_42 [425]);
assign l_41[394]    = ( l_42 [426]);
assign l_41[395]    = ( l_42 [427]);
assign l_41[396]    = ( l_42 [428]);
assign l_41[397]    = ( l_42 [429]);
assign l_41[398]    = ( l_42 [430]);
assign l_41[399]    = ( l_42 [431]);
assign l_41[400]    = ( l_42 [432]);
assign l_41[401]    = ( l_42 [433]);
assign l_41[402]    = ( l_42 [434]);
assign l_41[403]    = ( l_42 [435]);
assign l_41[404]    = ( l_42 [436]);
assign l_41[405]    = ( l_42 [437]);
assign l_41[406]    = ( l_42 [438]);
assign l_41[407]    = ( l_42 [439]);
assign l_41[408]    = ( l_42 [440]);
assign l_41[409]    = ( l_42 [441]);
assign l_41[410]    = ( l_42 [442]);
assign l_41[411]    = ( l_42 [443]);
assign l_41[412]    = ( l_42 [444]);
assign l_41[413]    = ( l_42 [445]);
assign l_41[414]    = ( l_42 [446]);
assign l_41[415]    = ( l_42 [447]);
assign l_41[416]    = ( l_42 [448]);
assign l_41[417]    = ( l_42 [449]);
assign l_41[418]    = ( l_42 [450]);
assign l_41[419]    = ( l_42 [451]);
assign l_41[420]    = ( l_42 [452]);
assign l_41[421]    = ( l_42 [453]);
assign l_41[422]    = ( l_42 [454]);
assign l_41[423]    = ( l_42 [455]);
assign l_41[424]    = ( l_42 [456]);
assign l_41[425]    = ( l_42 [457]);
assign l_41[426]    = ( l_42 [458]);
assign l_41[427]    = ( l_42 [459]);
assign l_41[428]    = ( l_42 [460]);
assign l_41[429]    = ( l_42 [461]);
assign l_41[430]    = ( l_42 [462]);
assign l_41[431]    = ( l_42 [463]);
assign l_41[432]    = ( l_42 [464]);
assign l_41[433]    = ( l_42 [465]);
assign l_41[434]    = ( l_42 [466]);
assign l_41[435]    = ( l_42 [467]);
assign l_41[436]    = ( l_42 [468]);
assign l_41[437]    = ( l_42 [469]);
assign l_41[438]    = ( l_42 [470]);
assign l_41[439]    = ( l_42 [471]);
assign l_41[440]    = ( l_42 [472]);
assign l_41[441]    = ( l_42 [473]);
assign l_41[442]    = ( l_42 [474]);
assign l_41[443]    = ( l_42 [475]);
assign l_41[444]    = ( l_42 [476]);
assign l_41[445]    = ( l_42 [477]);
assign l_41[446]    = ( l_42 [478]);
assign l_41[447]    = ( l_42 [479]);
assign l_41[448]    = ( l_42 [480]);
assign l_41[449]    = ( l_42 [481]);
assign l_41[450]    = ( l_42 [482]);
assign l_41[451]    = ( l_42 [483]);
assign l_41[452]    = ( l_42 [484]);
assign l_41[453]    = ( l_42 [485]);
assign l_41[454]    = ( l_42 [486]);
assign l_41[455]    = ( l_42 [487]);
assign l_41[456]    = ( l_42 [488]);
assign l_41[457]    = ( l_42 [489]);
assign l_41[458]    = ( l_42 [490]);
assign l_41[459]    = ( l_42 [491]);
assign l_41[460]    = ( l_42 [492]);
assign l_41[461]    = ( l_42 [493]);
assign l_41[462]    = ( l_42 [494]);
assign l_41[463]    = ( l_42 [495]);
assign l_41[464]    = ( l_42 [496]);
assign l_41[465]    = ( l_42 [497]);
assign l_41[466]    = ( l_42 [498]);
assign l_41[467]    = ( l_42 [499]);
assign l_41[468]    = ( l_42 [500]);
assign l_41[469]    = ( l_42 [501]);
assign l_41[470]    = ( l_42 [502]);
assign l_41[471]    = ( l_42 [503]);
assign l_41[472]    = ( l_42 [504]);
assign l_41[473]    = ( l_42 [505]);
assign l_41[474]    = ( l_42 [506]);
assign l_41[475]    = ( l_42 [507]);
assign l_41[476]    = ( l_42 [508]);
assign l_41[477]    = ( l_42 [509]);
assign l_41[478]    = ( l_42 [510]);
assign l_41[479]    = ( l_42 [511]);
assign l_41[480]    = ( l_42 [512]);
assign l_41[481]    = ( l_42 [513]);
assign l_41[482]    = ( l_42 [514]);
assign l_41[483]    = ( l_42 [515]);
assign l_41[484]    = ( l_42 [516]);
assign l_41[485]    = ( l_42 [517]);
assign l_41[486]    = ( l_42 [518]);
assign l_41[487]    = ( l_42 [519]);
assign l_41[488]    = ( l_42 [520]);
assign l_41[489]    = ( l_42 [521]);
assign l_41[490]    = ( l_42 [522]);
assign l_41[491]    = ( l_42 [523]);
assign l_41[492]    = ( l_42 [524]);
assign l_41[493]    = ( l_42 [525]);
assign l_41[494]    = ( l_42 [526]);
assign l_41[495]    = ( l_42 [527]);
assign l_41[496]    = ( l_42 [528]);
assign l_41[497]    = ( l_42 [529]);
assign l_41[498]    = ( l_42 [530]);
assign l_41[499]    = ( l_42 [531]);
assign l_41[500]    = ( l_42 [532]);
assign l_41[501]    = ( l_42 [533]);
assign l_41[502]    = ( l_42 [534]);
assign l_41[503]    = ( l_42 [535]);
assign l_41[504]    = ( l_42 [536]);
assign l_41[505]    = ( l_42 [537]);
assign l_41[506]    = ( l_42 [538]);
assign l_41[507]    = ( l_42 [539]);
assign l_41[508]    = ( l_42 [540]);
assign l_41[509]    = ( l_42 [541]);
assign l_41[510]    = ( l_42 [542]);
assign l_41[511]    = ( l_42 [543]);
assign l_41[512]    = ( l_42 [544]);
assign l_41[513]    = ( l_42 [545]);
assign l_41[514]    = ( l_42 [546]);
assign l_41[515]    = ( l_42 [547]);
assign l_41[516]    = ( l_42 [548]);
assign l_41[517]    = ( l_42 [549]);
assign l_41[518]    = ( l_42 [550]);
assign l_41[519]    = ( l_42 [551]);
assign l_41[520]    = ( l_42 [552]);
assign l_41[521]    = ( l_42 [553]);
assign l_41[522]    = ( l_42 [554]);
assign l_41[523]    = ( l_42 [555]);
assign l_41[524]    = ( l_42 [556]);
assign l_41[525]    = ( l_42 [557]);
assign l_41[526]    = ( l_42 [558]);
assign l_41[527]    = ( l_42 [559]);
assign l_41[528]    = ( l_42 [560]);
assign l_41[529]    = ( l_42 [561]);
assign l_41[530]    = ( l_42 [562]);
assign l_41[531]    = ( l_42 [563]);
assign l_41[532]    = ( l_42 [564]);
assign l_41[533]    = ( l_42 [565]);
assign l_41[534]    = ( l_42 [566]);
assign l_41[535]    = ( l_42 [567]);
assign l_41[536]    = ( l_42 [568]);
assign l_41[537]    = ( l_42 [569]);
assign l_41[538]    = ( l_42 [570]);
assign l_41[539]    = ( l_42 [571]);
assign l_41[540]    = ( l_42 [572]);
assign l_41[541]    = ( l_42 [573]);
assign l_41[542]    = ( l_42 [574]);
assign l_41[543]    = ( l_42 [575]);
assign l_41[544]    = ( l_42 [576]);
assign l_41[545]    = ( l_42 [577]);
assign l_41[546]    = ( l_42 [578]);
assign l_41[547]    = ( l_42 [579]);
assign l_41[548]    = ( l_42 [580]);
assign l_41[549]    = ( l_42 [581]);
assign l_41[550]    = ( l_42 [582]);
assign l_41[551]    = ( l_42 [583]);
assign l_41[552]    = ( l_42 [584]);
assign l_41[553]    = ( l_42 [585]);
assign l_41[554]    = ( l_42 [586]);
assign l_41[555]    = ( l_42 [587]);
assign l_41[556]    = ( l_42 [588]);
assign l_41[557]    = ( l_42 [589]);
assign l_41[558]    = ( l_42 [590]);
assign l_41[559]    = ( l_42 [591]);
assign l_41[560]    = ( l_42 [592]);
assign l_41[561]    = ( l_42 [593]);
assign l_41[562]    = ( l_42 [594]);
assign l_41[563]    = ( l_42 [595]);
assign l_41[564]    = ( l_42 [596]);
assign l_41[565]    = ( l_42 [597]);
assign l_41[566]    = ( l_42 [598]);
assign l_41[567]    = ( l_42 [599]);
assign l_41[568]    = ( l_42 [600]);
assign l_41[569]    = ( l_42 [601]);
assign l_41[570]    = ( l_42 [602]);
assign l_41[571]    = ( l_42 [603]);
assign l_41[572]    = ( l_42 [604]);
assign l_41[573]    = ( l_42 [605]);
assign l_41[574]    = ( l_42 [606]);
assign l_41[575]    = ( l_42 [607]);
assign l_41[576]    = ( l_42 [608]);
assign l_41[577]    = ( l_42 [609]);
assign l_41[578]    = ( l_42 [610]);
assign l_41[579]    = ( l_42 [611]);
assign l_41[580]    = ( l_42 [612]);
assign l_41[581]    = ( l_42 [613]);
assign l_41[582]    = ( l_42 [614]);
assign l_41[583]    = ( l_42 [615]);
assign l_41[584]    = ( l_42 [616]);
assign l_41[585]    = ( l_42 [617]);
assign l_41[586]    = ( l_42 [618]);
assign l_41[587]    = ( l_42 [619]);
assign l_41[588]    = ( l_42 [620]);
assign l_41[589]    = ( l_42 [621]);
assign l_41[590]    = ( l_42 [622]);
assign l_41[591]    = ( l_42 [623]);
assign l_41[592]    = ( l_42 [624]);
assign l_41[593]    = ( l_42 [625]);
assign l_41[594]    = ( l_42 [626]);
assign l_41[595]    = ( l_42 [627]);
assign l_41[596]    = ( l_42 [628]);
assign l_41[597]    = ( l_42 [629]);
assign l_41[598]    = ( l_42 [630]);
assign l_41[599]    = ( l_42 [631]);
assign l_41[600]    = ( l_42 [632]);
assign l_41[601]    = ( l_42 [633]);
assign l_41[602]    = ( l_42 [634]);
assign l_41[603]    = ( l_42 [635]);
assign l_41[604]    = ( l_42 [636]);
assign l_41[605]    = ( l_42 [637]);
assign l_41[606]    = ( l_42 [638]);
assign l_41[607]    = ( l_42 [639]);
assign l_41[608]    = ( l_42 [640]);
assign l_41[609]    = ( l_42 [641]);
assign l_41[610]    = ( l_42 [642]);
assign l_41[611]    = ( l_42 [643]);
assign l_41[612]    = ( l_42 [644]);
assign l_41[613]    = ( l_42 [645]);
assign l_41[614]    = ( l_42 [646]);
assign l_41[615]    = ( l_42 [647]);
assign l_41[616]    = ( l_42 [648]);
assign l_41[617]    = ( l_42 [649]);
assign l_41[618]    = ( l_42 [650]);
assign l_41[619]    = ( l_42 [651]);
assign l_41[620]    = ( l_42 [652]);
assign l_41[621]    = ( l_42 [653]);
assign l_41[622]    = ( l_42 [654]);
assign l_41[623]    = ( l_42 [655]);
assign l_41[624]    = ( l_42 [656]);
assign l_41[625]    = ( l_42 [657]);
assign l_41[626]    = ( l_42 [658]);
assign l_41[627]    = ( l_42 [659]);
assign l_41[628]    = ( l_42 [660]);
assign l_41[629]    = ( l_42 [661]);
assign l_41[630]    = ( l_42 [662]);
assign l_41[631]    = ( l_42 [663]);
assign l_41[632]    = ( l_42 [664]);
assign l_41[633]    = ( l_42 [665]);
assign l_41[634]    = ( l_42 [666]);
assign l_41[635]    = ( l_42 [667]);
assign l_41[636]    = ( l_42 [668]);
assign l_41[637]    = ( l_42 [669]);
assign l_41[638]    = ( l_42 [670]);
assign l_41[639]    = ( l_42 [671]);
assign l_41[640]    = ( l_42 [672]);
assign l_41[641]    = ( l_42 [673]);
assign l_41[642]    = ( l_42 [674]);
assign l_41[643]    = ( l_42 [675]);
assign l_41[644]    = ( l_42 [676]);
assign l_41[645]    = ( l_42 [677]);
assign l_41[646]    = ( l_42 [678]);
assign l_41[647]    = ( l_42 [679]);
assign l_41[648]    = ( l_42 [680]);
assign l_41[649]    = ( l_42 [681]);
assign l_41[650]    = ( l_42 [682]);
assign l_41[651]    = ( l_42 [683]);
assign l_41[652]    = ( l_42 [684]);
assign l_41[653]    = ( l_42 [685]);
assign l_41[654]    = ( l_42 [686]);
assign l_41[655]    = ( l_42 [687]);
assign l_41[656]    = ( l_42 [688]);
assign l_41[657]    = ( l_42 [689]);
assign l_41[658]    = ( l_42 [690]);
assign l_41[659]    = ( l_42 [691]);
assign l_41[660]    = ( l_42 [692]);
assign l_41[661]    = ( l_42 [693]);
assign l_41[662]    = ( l_42 [694]);
assign l_41[663]    = ( l_42 [695]);
assign l_41[664]    = ( l_42 [696]);
assign l_41[665]    = ( l_42 [697]);
assign l_41[666]    = ( l_42 [698]);
assign l_41[667]    = ( l_42 [699]);
assign l_41[668]    = ( l_42 [700]);
assign l_41[669]    = ( l_42 [701]);
assign l_41[670]    = ( l_42 [702]);
assign l_41[671]    = ( l_42 [703]);
assign l_41[672]    = ( l_42 [704]);
assign l_41[673]    = ( l_42 [705]);
assign l_41[674]    = ( l_42 [706]);
assign l_41[675]    = ( l_42 [707]);
assign l_41[676]    = ( l_42 [708]);
assign l_41[677]    = ( l_42 [709]);
assign l_41[678]    = ( l_42 [710]);
assign l_41[679]    = ( l_42 [711]);
assign l_41[680]    = ( l_42 [712]);
assign l_41[681]    = ( l_42 [713]);
assign l_41[682]    = ( l_42 [714]);
assign l_41[683]    = ( l_42 [715]);
assign l_41[684]    = ( l_42 [716]);
assign l_41[685]    = ( l_42 [717]);
assign l_41[686]    = ( l_42 [718]);
assign l_41[687]    = ( l_42 [719]);
assign l_41[688]    = ( l_42 [720]);
assign l_41[689]    = ( l_42 [721]);
assign l_41[690]    = ( l_42 [722]);
assign l_41[691]    = ( l_42 [723]);
assign l_41[692]    = ( l_42 [724]);
assign l_41[693]    = ( l_42 [725]);
assign l_41[694]    = ( l_42 [726]);
assign l_41[695]    = ( l_42 [727]);
assign l_41[696]    = ( l_42 [728]);
assign l_41[697]    = ( l_42 [729]);
assign l_41[698]    = ( l_42 [730]);
assign l_41[699]    = ( l_42 [731]);
assign l_41[700]    = ( l_42 [732]);
assign l_41[701]    = ( l_42 [733]);
assign l_41[702]    = ( l_42 [734]);
assign l_41[703]    = ( l_42 [735]);
assign l_41[704]    = ( l_42 [736]);
assign l_41[705]    = ( l_42 [737]);
assign l_41[706]    = ( l_42 [738]);
assign l_41[707]    = ( l_42 [739]);
assign l_41[708]    = ( l_42 [740]);
assign l_41[709]    = ( l_42 [741]);
assign l_41[710]    = ( l_42 [742]);
assign l_41[711]    = ( l_42 [743]);
assign l_41[712]    = ( l_42 [744]);
assign l_41[713]    = ( l_42 [745]);
assign l_41[714]    = ( l_42 [746]);
assign l_41[715]    = ( l_42 [747]);
assign l_41[716]    = ( l_42 [748]);
assign l_41[717]    = ( l_42 [749]);
assign l_41[718]    = ( l_42 [750]);
assign l_41[719]    = ( l_42 [751]);
assign l_41[720]    = ( l_42 [752]);
assign l_41[721]    = ( l_42 [753]);
assign l_41[722]    = ( l_42 [754]);
assign l_41[723]    = ( l_42 [755]);
assign l_41[724]    = ( l_42 [756]);
assign l_41[725]    = ( l_42 [757]);
assign l_41[726]    = ( l_42 [758]);
assign l_41[727]    = ( l_42 [759]);
assign l_41[728]    = ( l_42 [760]);
assign l_41[729]    = ( l_42 [761]);
assign l_41[730]    = ( l_42 [762]);
assign l_41[731]    = ( l_42 [763]);
assign l_41[732]    = ( l_42 [764]);
assign l_41[733]    = ( l_42 [765]);
assign l_41[734]    = ( l_42 [766]);
assign l_41[735]    = ( l_42 [767]);
assign l_41[736]    = ( l_42 [768]);
assign l_41[737]    = ( l_42 [769]);
assign l_41[738]    = ( l_42 [770]);
assign l_41[739]    = ( l_42 [771]);
assign l_41[740]    = ( l_42 [772]);
assign l_41[741]    = ( l_42 [773]);
assign l_41[742]    = ( l_42 [774]);
assign l_41[743]    = ( l_42 [775]);
assign l_41[744]    = ( l_42 [776]);
assign l_41[745]    = ( l_42 [777]);
assign l_41[746]    = ( l_42 [778]);
assign l_41[747]    = ( l_42 [779]);
assign l_41[748]    = ( l_42 [780]);
assign l_41[749]    = ( l_42 [781]);
assign l_41[750]    = ( l_42 [782]);
assign l_41[751]    = ( l_42 [783]);
assign l_41[752]    = ( l_42 [784]);
assign l_41[753]    = ( l_42 [785]);
assign l_41[754]    = ( l_42 [786]);
assign l_41[755]    = ( l_42 [787]);
assign l_41[756]    = ( l_42 [788]);
assign l_41[757]    = ( l_42 [789]);
assign l_41[758]    = ( l_42 [790]);
assign l_41[759]    = ( l_42 [791]);
assign l_41[760]    = ( l_42 [792]);
assign l_41[761]    = ( l_42 [793]);
assign l_41[762]    = ( l_42 [794]);
assign l_41[763]    = ( l_42 [795]);
assign l_41[764]    = ( l_42 [796]);
assign l_41[765]    = ( l_42 [797]);
assign l_41[766]    = ( l_42 [798]);
assign l_41[767]    = ( l_42 [799]);
assign l_41[768]    = ( l_42 [800]);
assign l_41[769]    = ( l_42 [801]);
assign l_41[770]    = ( l_42 [802]);
assign l_41[771]    = ( l_42 [803]);
assign l_41[772]    = ( l_42 [804]);
assign l_41[773]    = ( l_42 [805]);
assign l_41[774]    = ( l_42 [806]);
assign l_41[775]    = ( l_42 [807]);
assign l_41[776]    = ( l_42 [808]);
assign l_41[777]    = ( l_42 [809]);
assign l_41[778]    = ( l_42 [810]);
assign l_41[779]    = ( l_42 [811]);
assign l_41[780]    = ( l_42 [812]);
assign l_41[781]    = ( l_42 [813]);
assign l_41[782]    = ( l_42 [814]);
assign l_41[783]    = ( l_42 [815]);
assign l_41[784]    = ( l_42 [816]);
assign l_41[785]    = ( l_42 [817]);
assign l_41[786]    = ( l_42 [818]);
assign l_41[787]    = ( l_42 [819]);
assign l_41[788]    = ( l_42 [820]);
assign l_41[789]    = ( l_42 [821]);
assign l_41[790]    = ( l_42 [822]);
assign l_41[791]    = ( l_42 [823]);
assign l_41[792]    = ( l_42 [824]);
assign l_41[793]    = ( l_42 [825]);
assign l_41[794]    = ( l_42 [826]);
assign l_41[795]    = ( l_42 [827]);
assign l_41[796]    = ( l_42 [828]);
assign l_41[797]    = ( l_42 [829]);
assign l_41[798]    = ( l_42 [830]);
assign l_41[799]    = ( l_42 [831]);
assign l_41[800]    = ( l_42 [832]);
assign l_41[801]    = ( l_42 [833]);
assign l_41[802]    = ( l_42 [834]);
assign l_41[803]    = ( l_42 [835]);
assign l_41[804]    = ( l_42 [836]);
assign l_41[805]    = ( l_42 [837]);
assign l_41[806]    = ( l_42 [838]);
assign l_41[807]    = ( l_42 [839]);
assign l_41[808]    = ( l_42 [840]);
assign l_41[809]    = ( l_42 [841]);
assign l_41[810]    = ( l_42 [842]);
assign l_41[811]    = ( l_42 [843]);
assign l_41[812]    = ( l_42 [844]);
assign l_41[813]    = ( l_42 [845]);
assign l_41[814]    = ( l_42 [846]);
assign l_41[815]    = ( l_42 [847]);
assign l_41[816]    = ( l_42 [848]);
assign l_41[817]    = ( l_42 [849]);
assign l_41[818]    = ( l_42 [850]);
assign l_41[819]    = ( l_42 [851]);
assign l_41[820]    = ( l_42 [852]);
assign l_41[821]    = ( l_42 [853]);
assign l_41[822]    = ( l_42 [854]);
assign l_41[823]    = ( l_42 [855]);
assign l_41[824]    = ( l_42 [856]);
assign l_41[825]    = ( l_42 [857]);
assign l_41[826]    = ( l_42 [858]);
assign l_41[827]    = ( l_42 [859]);
assign l_41[828]    = ( l_42 [860]);
assign l_41[829]    = ( l_42 [861]);
assign l_41[830]    = ( l_42 [862]);
assign l_41[831]    = ( l_42 [863]);
assign l_41[832]    = ( l_42 [864]);
assign l_41[833]    = ( l_42 [865]);
assign l_41[834]    = ( l_42 [866]);
assign l_41[835]    = ( l_42 [867]);
assign l_41[836]    = ( l_42 [868]);
assign l_41[837]    = ( l_42 [869]);
assign l_41[838]    = ( l_42 [870]);
assign l_41[839]    = ( l_42 [871]);
assign l_41[840]    = ( l_42 [872]);
assign l_41[841]    = ( l_42 [873]);
assign l_41[842]    = ( l_42 [874]);
assign l_41[843]    = ( l_42 [875]);
assign l_41[844]    = ( l_42 [876]);
assign l_41[845]    = ( l_42 [877]);
assign l_41[846]    = ( l_42 [878]);
assign l_41[847]    = ( l_42 [879]);
assign l_41[848]    = ( l_42 [880]);
assign l_41[849]    = ( l_42 [881]);
assign l_41[850]    = ( l_42 [882]);
assign l_41[851]    = ( l_42 [883]);
assign l_41[852]    = ( l_42 [884]);
assign l_41[853]    = ( l_42 [885]);
assign l_41[854]    = ( l_42 [886]);
assign l_41[855]    = ( l_42 [887]);
assign l_41[856]    = ( l_42 [888]);
assign l_41[857]    = ( l_42 [889]);
assign l_41[858]    = ( l_42 [890]);
assign l_41[859]    = ( l_42 [891]);
assign l_41[860]    = ( l_42 [892]);
assign l_41[861]    = ( l_42 [893]);
assign l_41[862]    = ( l_42 [894]);
assign l_41[863]    = ( l_42 [895]);
assign l_41[864]    = ( l_42 [896]);
assign l_41[865]    = ( l_42 [897]);
assign l_41[866]    = ( l_42 [898]);
assign l_41[867]    = ( l_42 [899]);
assign l_41[868]    = ( l_42 [900]);
assign l_41[869]    = ( l_42 [901]);
assign l_41[870]    = ( l_42 [902]);
assign l_41[871]    = ( l_42 [903]);
assign l_41[872]    = ( l_42 [904]);
assign l_41[873]    = ( l_42 [905]);
assign l_41[874]    = ( l_42 [906]);
assign l_41[875]    = ( l_42 [907]);
assign l_41[876]    = ( l_42 [908]);
assign l_41[877]    = ( l_42 [909]);
assign l_41[878]    = ( l_42 [910]);
assign l_41[879]    = ( l_42 [911]);
assign l_41[880]    = ( l_42 [912]);
assign l_41[881]    = ( l_42 [913]);
assign l_41[882]    = ( l_42 [914]);
assign l_41[883]    = ( l_42 [915]);
assign l_41[884]    = ( l_42 [916]);
assign l_41[885]    = ( l_42 [917]);
assign l_41[886]    = ( l_42 [918]);
assign l_41[887]    = ( l_42 [919]);
assign l_41[888]    = ( l_42 [920]);
assign l_41[889]    = ( l_42 [921]);
assign l_41[890]    = ( l_42 [922]);
assign l_41[891]    = ( l_42 [923]);
assign l_41[892]    = ( l_42 [924]);
assign l_41[893]    = ( l_42 [925]);
assign l_41[894]    = ( l_42 [926]);
assign l_41[895]    = ( l_42 [927]);
assign l_41[896]    = ( l_42 [928]);
assign l_41[897]    = ( l_42 [929]);
assign l_41[898]    = ( l_42 [930]);
assign l_41[899]    = ( l_42 [931]);
assign l_41[900]    = ( l_42 [932]);
assign l_41[901]    = ( l_42 [933]);
assign l_41[902]    = ( l_42 [934]);
assign l_41[903]    = ( l_42 [935]);
assign l_41[904]    = ( l_42 [936]);
assign l_41[905]    = ( l_42 [937]);
assign l_41[906]    = ( l_42 [938]);
assign l_41[907]    = ( l_42 [939]);
assign l_41[908]    = ( l_42 [940]);
assign l_41[909]    = ( l_42 [941]);
assign l_41[910]    = ( l_42 [942]);
assign l_41[911]    = ( l_42 [943]);
assign l_41[912]    = ( l_42 [944]);
assign l_41[913]    = ( l_42 [945]);
assign l_41[914]    = ( l_42 [946]);
assign l_41[915]    = ( l_42 [947]);
assign l_41[916]    = ( l_42 [948]);
assign l_41[917]    = ( l_42 [949]);
assign l_41[918]    = ( l_42 [950]);
assign l_41[919]    = ( l_42 [951]);
assign l_41[920]    = ( l_42 [952]);
assign l_41[921]    = ( l_42 [953]);
assign l_41[922]    = ( l_42 [954]);
assign l_41[923]    = ( l_42 [955]);
assign l_41[924]    = ( l_42 [956]);
assign l_41[925]    = ( l_42 [957]);
assign l_41[926]    = ( l_42 [958]);
assign l_41[927]    = ( l_42 [959]);
assign l_41[928]    = ( l_42 [960]);
assign l_41[929]    = ( l_42 [961]);
assign l_41[930]    = ( l_42 [962]);
assign l_41[931]    = ( l_42 [963]);
assign l_41[932]    = ( l_42 [964]);
assign l_41[933]    = ( l_42 [965]);
assign l_41[934]    = ( l_42 [966]);
assign l_41[935]    = ( l_42 [967]);
assign l_41[936]    = ( l_42 [968]);
assign l_41[937]    = ( l_42 [969]);
assign l_41[938]    = ( l_42 [970]);
assign l_41[939]    = ( l_42 [971]);
assign l_41[940]    = ( l_42 [972]);
assign l_41[941]    = ( l_42 [973]);
assign l_41[942]    = ( l_42 [974]);
assign l_41[943]    = ( l_42 [975]);
assign l_41[944]    = ( l_42 [976]);
assign l_41[945]    = ( l_42 [977]);
assign l_41[946]    = ( l_42 [978]);
assign l_41[947]    = ( l_42 [979]);
assign l_41[948]    = ( l_42 [980]);
assign l_41[949]    = ( l_42 [981]);
assign l_41[950]    = ( l_42 [982]);
assign l_41[951]    = ( l_42 [983]);
assign l_41[952]    = ( l_42 [984]);
assign l_41[953]    = ( l_42 [985]);
assign l_41[954]    = ( l_42 [986]);
assign l_41[955]    = ( l_42 [987]);
assign l_41[956]    = ( l_42 [988]);
assign l_41[957]    = ( l_42 [989]);
assign l_41[958]    = ( l_42 [990]);
assign l_41[959]    = ( l_42 [991]);
assign l_41[960]    = ( l_42 [992]);
assign l_41[961]    = ( l_42 [993]);
assign l_41[962]    = ( l_42 [994]);
assign l_41[963]    = ( l_42 [995]);
assign l_41[964]    = ( l_42 [996]);
assign l_41[965]    = ( l_42 [997]);
assign l_41[966]    = ( l_42 [998]);
assign l_41[967]    = ( l_42 [999]);
assign l_41[968]    = ( l_42 [1000]);
assign l_41[969]    = ( l_42 [1001]);
assign l_41[970]    = ( l_42 [1002]);
assign l_41[971]    = ( l_42 [1003]);
assign l_41[972]    = ( l_42 [1004]);
assign l_41[973]    = ( l_42 [1005]);
assign l_41[974]    = ( l_42 [1006]);
assign l_41[975]    = ( l_42 [1007]);
assign l_41[976]    = ( l_42 [1008]);
assign l_41[977]    = ( l_42 [1009]);
assign l_41[978]    = ( l_42 [1010]);
assign l_41[979]    = ( l_42 [1011]);
assign l_41[980]    = ( l_42 [1012]);
assign l_41[981]    = ( l_42 [1013]);
assign l_41[982]    = ( l_42 [1014]);
assign l_41[983]    = ( l_42 [1015]);
assign l_41[984]    = ( l_42 [1016]);
assign l_41[985]    = ( l_42 [1017]);
assign l_41[986]    = ( l_42 [1018]);
assign l_41[987]    = ( l_42 [1019]);
assign l_41[988]    = ( l_42 [1020]);
assign l_41[989]    = ( l_42 [1021]);
assign l_41[990]    = ( l_42 [1022]);
assign l_41[991]    = ( l_42 [1023]);
assign l_41[992]    = ( l_42 [1024]);
assign l_41[993]    = ( l_42 [1025]);
assign l_41[994]    = ( l_42 [1026]);
assign l_41[995]    = ( l_42 [1027]);
assign l_41[996]    = ( l_42 [1028]);
assign l_41[997]    = ( l_42 [1029]);
assign l_41[998]    = ( l_42 [1030]);
assign l_41[999]    = ( l_42 [1031]);
assign l_41[1000]    = ( l_42 [1032]);
assign l_41[1001]    = ( l_42 [1033]);
assign l_41[1002]    = ( l_42 [1034]);
assign l_41[1003]    = ( l_42 [1035]);
assign l_41[1004]    = ( l_42 [1036]);
assign l_41[1005]    = ( l_42 [1037]);
assign l_41[1006]    = ( l_42 [1038]);
assign l_41[1007]    = ( l_42 [1039]);
assign l_41[1008]    = ( l_42 [1040]);
assign l_41[1009]    = ( l_42 [1041]);
assign l_41[1010]    = ( l_42 [1042]);
assign l_41[1011]    = ( l_42 [1043]);
assign l_41[1012]    = ( l_42 [1044]);
assign l_41[1013]    = ( l_42 [1045]);
assign l_41[1014]    = ( l_42 [1046]);
assign l_41[1015]    = ( l_42 [1047]);
assign l_41[1016]    = ( l_42 [1048]);
assign l_41[1017]    = ( l_42 [1049]);
assign l_41[1018]    = ( l_42 [1050]);
assign l_41[1019]    = ( l_42 [1051]);
assign l_41[1020]    = ( l_42 [1052]);
assign l_41[1021]    = ( l_42 [1053]);
assign l_41[1022]    = ( l_42 [1054]);
assign l_41[1023]    = ( l_42 [1055]);
assign l_41[1024]    = ( l_42 [1056]);
assign l_41[1025]    = ( l_42 [1057]);
assign l_41[1026]    = ( l_42 [1058]);
assign l_41[1027]    = ( l_42 [1059]);
assign l_41[1028]    = ( l_42 [1060]);
assign l_41[1029]    = ( l_42 [1061]);
assign l_41[1030]    = ( l_42 [1062]);
assign l_41[1031]    = ( l_42 [1063]);
assign l_41[1032]    = ( l_42 [1064]);
assign l_41[1033]    = ( l_42 [1065]);
assign l_41[1034]    = ( l_42 [1066]);
assign l_41[1035]    = ( l_42 [1067]);
assign l_41[1036]    = ( l_42 [1068]);
assign l_41[1037]    = ( l_42 [1069]);
assign l_41[1038]    = ( l_42 [1070]);
assign l_41[1039]    = ( l_42 [1071]);
assign l_41[1040]    = ( l_42 [1072]);
assign l_41[1041]    = ( l_42 [1073]);
assign l_41[1042]    = ( l_42 [1074]);
assign l_41[1043]    = ( l_42 [1075]);
assign l_41[1044]    = ( l_42 [1076]);
assign l_41[1045]    = ( l_42 [1077]);
assign l_41[1046]    = ( l_42 [1078]);
assign l_41[1047]    = ( l_42 [1079]);
assign l_41[1048]    = ( l_42 [1080]);
assign l_41[1049]    = ( l_42 [1081]);
assign l_41[1050]    = ( l_42 [1082]);
assign l_41[1051]    = ( l_42 [1083]);
assign l_41[1052]    = ( l_42 [1084]);
assign l_41[1053]    = ( l_42 [1085]);
assign l_41[1054]    = ( l_42 [1086]);
assign l_41[1055]    = ( l_42 [1087]);
assign l_41[1056]    = ( l_42 [1088]);
assign l_41[1057]    = ( l_42 [1089]);
assign l_41[1058]    = ( l_42 [1090]);
assign l_41[1059]    = ( l_42 [1091]);
assign l_41[1060]    = ( l_42 [1092]);
assign l_41[1061]    = ( l_42 [1093]);
assign l_41[1062]    = ( l_42 [1094]);
assign l_41[1063]    = ( l_42 [1095]);
assign l_41[1064]    = ( l_42 [1096]);
assign l_41[1065]    = ( l_42 [1097]);
assign l_41[1066]    = ( l_42 [1098]);
assign l_41[1067]    = ( l_42 [1099]);
assign l_41[1068]    = ( l_42 [1100]);
assign l_41[1069]    = ( l_42 [1101]);
assign l_41[1070]    = ( l_42 [1102]);
assign l_41[1071]    = ( l_42 [1103]);
assign l_41[1072]    = ( l_42 [1104]);
assign l_41[1073]    = ( l_42 [1105]);
assign l_41[1074]    = ( l_42 [1106]);
assign l_41[1075]    = ( l_42 [1107]);
assign l_41[1076]    = ( l_42 [1108]);
assign l_41[1077]    = ( l_42 [1109]);
assign l_41[1078]    = ( l_42 [1110]);
assign l_41[1079]    = ( l_42 [1111]);
assign l_41[1080]    = ( l_42 [1112]);
assign l_41[1081]    = ( l_42 [1113]);
assign l_41[1082]    = ( l_42 [1114]);
assign l_41[1083]    = ( l_42 [1115]);
assign l_41[1084]    = ( l_42 [1116]);
assign l_41[1085]    = ( l_42 [1117]);
assign l_41[1086]    = ( l_42 [1118]);
assign l_41[1087]    = ( l_42 [1119]);
assign l_41[1088]    = ( l_42 [1120]);
assign l_41[1089]    = ( l_42 [1121]);
assign l_41[1090]    = ( l_42 [1122]);
assign l_41[1091]    = ( l_42 [1123]);
assign l_41[1092]    = ( l_42 [1124]);
assign l_41[1093]    = ( l_42 [1125]);
assign l_41[1094]    = ( l_42 [1126]);
assign l_41[1095]    = ( l_42 [1127]);
assign l_41[1096]    = ( l_42 [1128]);
assign l_41[1097]    = ( l_42 [1129]);
assign l_41[1098]    = ( l_42 [1130]);
assign l_41[1099]    = ( l_42 [1131]);
assign l_41[1100]    = ( l_42 [1132]);
assign l_41[1101]    = ( l_42 [1133]);
assign l_41[1102]    = ( l_42 [1134]);
assign l_41[1103]    = ( l_42 [1135]);
assign l_41[1104]    = ( l_42 [1136]);
assign l_41[1105]    = ( l_42 [1137]);
assign l_41[1106]    = ( l_42 [1138]);
assign l_41[1107]    = ( l_42 [1139]);
assign l_41[1108]    = ( l_42 [1140]);
assign l_41[1109]    = ( l_42 [1141]);
assign l_41[1110]    = ( l_42 [1142]);
assign l_41[1111]    = ( l_42 [1143]);
assign l_41[1112]    = ( l_42 [1144]);
assign l_41[1113]    = ( l_42 [1145]);
assign l_41[1114]    = ( l_42 [1146]);
assign l_41[1115]    = ( l_42 [1147]);
assign l_41[1116]    = ( l_42 [1148]);
assign l_41[1117]    = ( l_42 [1149]);
assign l_41[1118]    = ( l_42 [1150]);
assign l_41[1119]    = ( l_42 [1151]);
assign l_41[1120]    = ( l_42 [1152]);
assign l_41[1121]    = ( l_42 [1153]);
assign l_41[1122]    = ( l_42 [1154]);
assign l_41[1123]    = ( l_42 [1155]);
assign l_41[1124]    = ( l_42 [1156]);
assign l_41[1125]    = ( l_42 [1157]);
assign l_41[1126]    = ( l_42 [1158]);
assign l_41[1127]    = ( l_42 [1159]);
assign l_41[1128]    = ( l_42 [1160]);
assign l_41[1129]    = ( l_42 [1161]);
assign l_41[1130]    = ( l_42 [1162]);
assign l_41[1131]    = ( l_42 [1163]);
assign l_41[1132]    = ( l_42 [1164]);
assign l_41[1133]    = ( l_42 [1165]);
assign l_41[1134]    = ( l_42 [1166]);
assign l_41[1135]    = ( l_42 [1167]);
assign l_41[1136]    = ( l_42 [1168]);
assign l_41[1137]    = ( l_42 [1169]);
assign l_41[1138]    = ( l_42 [1170]);
assign l_41[1139]    = ( l_42 [1171]);
assign l_41[1140]    = ( l_42 [1172]);
assign l_41[1141]    = ( l_42 [1173]);
assign l_41[1142]    = ( l_42 [1174]);
assign l_41[1143]    = ( l_42 [1175]);
assign l_41[1144]    = ( l_42 [1176]);
assign l_41[1145]    = ( l_42 [1177]);
assign l_41[1146]    = ( l_42 [1178]);
assign l_41[1147]    = ( l_42 [1179]);
assign l_41[1148]    = ( l_42 [1180]);
assign l_41[1149]    = ( l_42 [1181]);
assign l_41[1150]    = ( l_42 [1182]);
assign l_41[1151]    = ( l_42 [1183]);
assign l_41[1152]    = ( l_42 [1184]);
assign l_41[1153]    = ( l_42 [1185]);
assign l_41[1154]    = ( l_42 [1186]);
assign l_41[1155]    = ( l_42 [1187]);
assign l_41[1156]    = ( l_42 [1188]);
assign l_41[1157]    = ( l_42 [1189]);
assign l_41[1158]    = ( l_42 [1190]);
assign l_41[1159]    = ( l_42 [1191]);
assign l_41[1160]    = ( l_42 [1192]);
assign l_41[1161]    = ( l_42 [1193]);
assign l_41[1162]    = ( l_42 [1194]);
assign l_41[1163]    = ( l_42 [1195]);
assign l_41[1164]    = ( l_42 [1196]);
assign l_41[1165]    = ( l_42 [1197]);
assign l_41[1166]    = ( l_42 [1198]);
assign l_41[1167]    = ( l_42 [1199]);
assign l_41[1168]    = ( l_42 [1200]);
assign l_41[1169]    = ( l_42 [1201]);
assign l_41[1170]    = ( l_42 [1202]);
assign l_41[1171]    = ( l_42 [1203]);
assign l_41[1172]    = ( l_42 [1204]);
assign l_41[1173]    = ( l_42 [1205]);
assign l_41[1174]    = ( l_42 [1206]);
assign l_41[1175]    = ( l_42 [1207]);
assign l_41[1176]    = ( l_42 [1208]);
assign l_41[1177]    = ( l_42 [1209]);
assign l_41[1178]    = ( l_42 [1210]);
assign l_41[1179]    = ( l_42 [1211]);
assign l_41[1180]    = ( l_42 [1212]);
assign l_41[1181]    = ( l_42 [1213]);
assign l_41[1182]    = ( l_42 [1214]);
assign l_41[1183]    = ( l_42 [1215]);
assign l_41[1184]    = ( l_42 [1216]);
assign l_41[1185]    = ( l_42 [1217]);
assign l_41[1186]    = ( l_42 [1218]);
assign l_41[1187]    = ( l_42 [1219]);
assign l_41[1188]    = ( l_42 [1220]);
assign l_41[1189]    = ( l_42 [1221]);
assign l_41[1190]    = ( l_42 [1222]);
assign l_41[1191]    = ( l_42 [1223]);
assign l_41[1192]    = ( l_42 [1224]);
assign l_41[1193]    = ( l_42 [1225]);
assign l_41[1194]    = ( l_42 [1226]);
assign l_41[1195]    = ( l_42 [1227]);
assign l_41[1196]    = ( l_42 [1228]);
assign l_41[1197]    = ( l_42 [1229]);
assign l_41[1198]    = ( l_42 [1230]);
assign l_41[1199]    = ( l_42 [1231]);
assign l_41[1200]    = ( l_42 [1232]);
assign l_41[1201]    = ( l_42 [1233]);
assign l_41[1202]    = ( l_42 [1234]);
assign l_41[1203]    = ( l_42 [1235]);
assign l_41[1204]    = ( l_42 [1236]);
assign l_41[1205]    = ( l_42 [1237]);
assign l_41[1206]    = ( l_42 [1238]);
assign l_41[1207]    = ( l_42 [1239]);
assign l_41[1208]    = ( l_42 [1240]);
assign l_41[1209]    = ( l_42 [1241]);
assign l_41[1210]    = ( l_42 [1242]);
assign l_41[1211]    = ( l_42 [1243]);
assign l_41[1212]    = ( l_42 [1244]);
assign l_41[1213]    = ( l_42 [1245]);
assign l_41[1214]    = ( l_42 [1246]);
assign l_41[1215]    = ( l_42 [1247]);
assign l_41[1216]    = ( l_42 [1248]);
assign l_41[1217]    = ( l_42 [1249]);
assign l_41[1218]    = ( l_42 [1250]);
assign l_41[1219]    = ( l_42 [1251]);
assign l_41[1220]    = ( l_42 [1252]);
assign l_41[1221]    = ( l_42 [1253]);
assign l_41[1222]    = ( l_42 [1254]);
assign l_41[1223]    = ( l_42 [1255]);
assign l_41[1224]    = ( l_42 [1256]);
assign l_41[1225]    = ( l_42 [1257]);
assign l_41[1226]    = ( l_42 [1258]);
assign l_41[1227]    = ( l_42 [1259]);
assign l_41[1228]    = ( l_42 [1260]);
assign l_41[1229]    = ( l_42 [1261]);
assign l_41[1230]    = ( l_42 [1262]);
assign l_41[1231]    = ( l_42 [1263]);
assign l_41[1232]    = ( l_42 [1264]);
assign l_41[1233]    = ( l_42 [1265]);
assign l_41[1234]    = ( l_42 [1266]);
assign l_41[1235]    = ( l_42 [1267]);
assign l_41[1236]    = ( l_42 [1268]);
assign l_41[1237]    = ( l_42 [1269]);
assign l_41[1238]    = ( l_42 [1270]);
assign l_41[1239]    = ( l_42 [1271]);
assign l_41[1240]    = ( l_42 [1272]);
assign l_41[1241]    = ( l_42 [1273]);
assign l_41[1242]    = ( l_42 [1274]);
assign l_41[1243]    = ( l_42 [1275]);
assign l_41[1244]    = ( l_42 [1276]);
assign l_41[1245]    = ( l_42 [1277]);
assign l_41[1246]    = ( l_42 [1278]);
assign l_41[1247]    = ( l_42 [1279]);
assign l_41[1248]    = ( l_42 [1280]);
assign l_41[1249]    = ( l_42 [1281]);
assign l_41[1250]    = ( l_42 [1282]);
assign l_41[1251]    = ( l_42 [1283]);
assign l_41[1252]    = ( l_42 [1284]);
assign l_41[1253]    = ( l_42 [1285]);
assign l_41[1254]    = ( l_42 [1286]);
assign l_41[1255]    = ( l_42 [1287]);
assign l_41[1256]    = ( l_42 [1288]);
assign l_41[1257]    = ( l_42 [1289]);
assign l_41[1258]    = ( l_42 [1290]);
assign l_41[1259]    = ( l_42 [1291]);
assign l_41[1260]    = ( l_42 [1292]);
assign l_41[1261]    = ( l_42 [1293]);
assign l_41[1262]    = ( l_42 [1294]);
assign l_41[1263]    = ( l_42 [1295]);
assign l_41[1264]    = ( l_42 [1296]);
assign l_41[1265]    = ( l_42 [1297]);
assign l_41[1266]    = ( l_42 [1298]);
assign l_41[1267]    = ( l_42 [1299]);
assign l_41[1268]    = ( l_42 [1300]);
assign l_41[1269]    = ( l_42 [1301]);
assign l_41[1270]    = ( l_42 [1302]);
assign l_41[1271]    = ( l_42 [1303]);
assign l_41[1272]    = ( l_42 [1304]);
assign l_41[1273]    = ( l_42 [1305]);
assign l_41[1274]    = ( l_42 [1306]);
assign l_41[1275]    = ( l_42 [1307]);
assign l_41[1276]    = ( l_42 [1308]);
assign l_41[1277]    = ( l_42 [1309]);
assign l_41[1278]    = ( l_42 [1310]);
assign l_41[1279]    = ( l_42 [1311]);
assign l_41[1280]    = ( l_42 [1312]);
assign l_41[1281]    = ( l_42 [1313]);
assign l_41[1282]    = ( l_42 [1314]);
assign l_41[1283]    = ( l_42 [1315]);
assign l_41[1284]    = ( l_42 [1316]);
assign l_41[1285]    = ( l_42 [1317]);
assign l_41[1286]    = ( l_42 [1318]);
assign l_41[1287]    = ( l_42 [1319]);
assign l_41[1288]    = ( l_42 [1320]);
assign l_41[1289]    = ( l_42 [1321]);
assign l_41[1290]    = ( l_42 [1322]);
assign l_41[1291]    = ( l_42 [1323]);
assign l_41[1292]    = ( l_42 [1324]);
assign l_41[1293]    = ( l_42 [1325]);
assign l_41[1294]    = ( l_42 [1326]);
assign l_41[1295]    = ( l_42 [1327]);
assign l_41[1296]    = ( l_42 [1328]);
assign l_41[1297]    = ( l_42 [1329]);
assign l_41[1298]    = ( l_42 [1330]);
assign l_41[1299]    = ( l_42 [1331]);
assign l_41[1300]    = ( l_42 [1332]);
assign l_41[1301]    = ( l_42 [1333]);
assign l_41[1302]    = ( l_42 [1334]);
assign l_41[1303]    = ( l_42 [1335]);
assign l_41[1304]    = ( l_42 [1336]);
assign l_41[1305]    = ( l_42 [1337]);
assign l_41[1306]    = ( l_42 [1338]);
assign l_41[1307]    = ( l_42 [1339]);
assign l_41[1308]    = ( l_42 [1340]);
assign l_41[1309]    = ( l_42 [1341]);
assign l_41[1310]    = ( l_42 [1342]);
assign l_41[1311]    = ( l_42 [1343]);
assign l_41[1312]    = ( l_42 [1344]);
assign l_41[1313]    = ( l_42 [1345]);
assign l_41[1314]    = ( l_42 [1346]);
assign l_41[1315]    = ( l_42 [1347]);
assign l_41[1316]    = ( l_42 [1348]);
assign l_41[1317]    = ( l_42 [1349]);
assign l_41[1318]    = ( l_42 [1350]);
assign l_41[1319]    = ( l_42 [1351]);
assign l_41[1320]    = ( l_42 [1352]);
assign l_41[1321]    = ( l_42 [1353]);
assign l_41[1322]    = ( l_42 [1354]);
assign l_41[1323]    = ( l_42 [1355]);
assign l_41[1324]    = ( l_42 [1356]);
assign l_41[1325]    = ( l_42 [1357]);
assign l_41[1326]    = ( l_42 [1358]);
assign l_41[1327]    = ( l_42 [1359]);
assign l_41[1328]    = ( l_42 [1360]);
assign l_41[1329]    = ( l_42 [1361]);
assign l_41[1330]    = ( l_42 [1362]);
assign l_41[1331]    = ( l_42 [1363]);
assign l_41[1332]    = ( l_42 [1364]);
assign l_41[1333]    = ( l_42 [1365]);
assign l_41[1334]    = ( l_42 [1366]);
assign l_41[1335]    = ( l_42 [1367]);
assign l_41[1336]    = ( l_42 [1368]);
assign l_41[1337]    = ( l_42 [1369]);
assign l_41[1338]    = ( l_42 [1370]);
assign l_41[1339]    = ( l_42 [1371]);
assign l_41[1340]    = ( l_42 [1372]);
assign l_41[1341]    = ( l_42 [1373]);
assign l_41[1342]    = ( l_42 [1374]);
assign l_41[1343]    = ( l_42 [1375]);
assign l_41[1344]    = ( l_42 [1376]);
assign l_41[1345]    = ( l_42 [1377]);
assign l_41[1346]    = ( l_42 [1378]);
assign l_41[1347]    = ( l_42 [1379]);
assign l_41[1348]    = ( l_42 [1380]);
assign l_41[1349]    = ( l_42 [1381]);
assign l_41[1350]    = ( l_42 [1382]);
assign l_41[1351]    = ( l_42 [1383]);
assign l_41[1352]    = ( l_42 [1384]);
assign l_41[1353]    = ( l_42 [1385]);
assign l_41[1354]    = ( l_42 [1386]);
assign l_41[1355]    = ( l_42 [1387]);
assign l_41[1356]    = ( l_42 [1388]);
assign l_41[1357]    = ( l_42 [1389]);
assign l_41[1358]    = ( l_42 [1390]);
assign l_41[1359]    = ( l_42 [1391]);
assign l_41[1360]    = ( l_42 [1392]);
assign l_41[1361]    = ( l_42 [1393]);
assign l_41[1362]    = ( l_42 [1394]);
assign l_41[1363]    = ( l_42 [1395]);
assign l_41[1364]    = ( l_42 [1396]);
assign l_41[1365]    = ( l_42 [1397]);
assign l_41[1366]    = ( l_42 [1398]);
assign l_41[1367]    = ( l_42 [1399]);
assign l_41[1368]    = ( l_42 [1400]);
assign l_41[1369]    = ( l_42 [1401]);
assign l_41[1370]    = ( l_42 [1402]);
assign l_41[1371]    = ( l_42 [1403]);
assign l_41[1372]    = ( l_42 [1404]);
assign l_41[1373]    = ( l_42 [1405]);
assign l_41[1374]    = ( l_42 [1406]);
assign l_41[1375]    = ( l_42 [1407]);
assign l_41[1376]    = ( l_42 [1408]);
assign l_41[1377]    = ( l_42 [1409]);
assign l_41[1378]    = ( l_42 [1410]);
assign l_41[1379]    = ( l_42 [1411]);
assign l_41[1380]    = ( l_42 [1412]);
assign l_41[1381]    = ( l_42 [1413]);
assign l_41[1382]    = ( l_42 [1414]);
assign l_41[1383]    = ( l_42 [1415]);
assign l_41[1384]    = ( l_42 [1416]);
assign l_41[1385]    = ( l_42 [1417]);
assign l_41[1386]    = ( l_42 [1418]);
assign l_41[1387]    = ( l_42 [1419]);
assign l_41[1388]    = ( l_42 [1420]);
assign l_41[1389]    = ( l_42 [1421]);
assign l_41[1390]    = ( l_42 [1422]);
assign l_41[1391]    = ( l_42 [1423]);
assign l_41[1392]    = ( l_42 [1424]);
assign l_41[1393]    = ( l_42 [1425]);
assign l_41[1394]    = ( l_42 [1426]);
assign l_41[1395]    = ( l_42 [1427]);
assign l_41[1396]    = ( l_42 [1428]);
assign l_41[1397]    = ( l_42 [1429]);
assign l_41[1398]    = ( l_42 [1430]);
assign l_41[1399]    = ( l_42 [1431]);
assign l_41[1400]    = ( l_42 [1432]);
assign l_41[1401]    = ( l_42 [1433]);
assign l_41[1402]    = ( l_42 [1434]);
assign l_41[1403]    = ( l_42 [1435]);
assign l_41[1404]    = ( l_42 [1436]);
assign l_41[1405]    = ( l_42 [1437]);
assign l_41[1406]    = ( l_42 [1438]);
assign l_41[1407]    = ( l_42 [1439]);
assign l_41[1408]    = ( l_42 [1440]);
assign l_41[1409]    = ( l_42 [1441]);
assign l_41[1410]    = ( l_42 [1442]);
assign l_41[1411]    = ( l_42 [1443]);
assign l_41[1412]    = ( l_42 [1444]);
assign l_41[1413]    = ( l_42 [1445]);
assign l_41[1414]    = ( l_42 [1446]);
assign l_41[1415]    = ( l_42 [1447]);
assign l_41[1416]    = ( l_42 [1448]);
assign l_41[1417]    = ( l_42 [1449]);
assign l_41[1418]    = ( l_42 [1450]);
assign l_41[1419]    = ( l_42 [1451]);
assign l_41[1420]    = ( l_42 [1452]);
assign l_41[1421]    = ( l_42 [1453]);
assign l_41[1422]    = ( l_42 [1454]);
assign l_41[1423]    = ( l_42 [1455]);
assign l_41[1424]    = ( l_42 [1456]);
assign l_41[1425]    = ( l_42 [1457]);
assign l_41[1426]    = ( l_42 [1458]);
assign l_41[1427]    = ( l_42 [1459]);
assign l_41[1428]    = ( l_42 [1460]);
assign l_41[1429]    = ( l_42 [1461]);
assign l_41[1430]    = ( l_42 [1462]);
assign l_41[1431]    = ( l_42 [1463]);
assign l_41[1432]    = ( l_42 [1464]);
assign l_41[1433]    = ( l_42 [1465]);
assign l_41[1434]    = ( l_42 [1466]);
assign l_41[1435]    = ( l_42 [1467]);
assign l_41[1436]    = ( l_42 [1468]);
assign l_41[1437]    = ( l_42 [1469]);
assign l_41[1438]    = ( l_42 [1470]);
assign l_41[1439]    = ( l_42 [1471]);
assign l_41[1440]    = ( l_42 [1472]);
assign l_41[1441]    = ( l_42 [1473]);
assign l_41[1442]    = ( l_42 [1474]);
assign l_41[1443]    = ( l_42 [1475]);
assign l_41[1444]    = ( l_42 [1476]);
assign l_41[1445]    = ( l_42 [1477]);
assign l_41[1446]    = ( l_42 [1478]);
assign l_41[1447]    = ( l_42 [1479]);
assign l_41[1448]    = ( l_42 [1480]);
assign l_41[1449]    = ( l_42 [1481]);
assign l_41[1450]    = ( l_42 [1482]);
assign l_41[1451]    = ( l_42 [1483]);
assign l_41[1452]    = ( l_42 [1484]);
assign l_41[1453]    = ( l_42 [1485]);
assign l_41[1454]    = ( l_42 [1486]);
assign l_41[1455]    = ( l_42 [1487]);
assign l_41[1456]    = ( l_42 [1488]);
assign l_41[1457]    = ( l_42 [1489]);
assign l_41[1458]    = ( l_42 [1490]);
assign l_41[1459]    = ( l_42 [1491]);
assign l_41[1460]    = ( l_42 [1492]);
assign l_41[1461]    = ( l_42 [1493]);
assign l_41[1462]    = ( l_42 [1494]);
assign l_41[1463]    = ( l_42 [1495]);
assign l_41[1464]    = ( l_42 [1496]);
assign l_41[1465]    = ( l_42 [1497]);
assign l_41[1466]    = ( l_42 [1498]);
assign l_41[1467]    = ( l_42 [1499]);
assign l_41[1468]    = ( l_42 [1500]);
assign l_41[1469]    = ( l_42 [1501]);
assign l_41[1470]    = ( l_42 [1502]);
assign l_41[1471]    = ( l_42 [1503]);
assign l_41[1472]    = ( l_42 [1504]);
assign l_41[1473]    = ( l_42 [1505]);
assign l_41[1474]    = ( l_42 [1506]);
assign l_41[1475]    = ( l_42 [1507]);
assign l_41[1476]    = ( l_42 [1508]);
assign l_41[1477]    = ( l_42 [1509]);
assign l_41[1478]    = ( l_42 [1510]);
assign l_41[1479]    = ( l_42 [1511]);
assign l_41[1480]    = ( l_42 [1512]);
assign l_41[1481]    = ( l_42 [1513]);
assign l_41[1482]    = ( l_42 [1514]);
assign l_41[1483]    = ( l_42 [1515]);
assign l_41[1484]    = ( l_42 [1516]);
assign l_41[1485]    = ( l_42 [1517]);
assign l_41[1486]    = ( l_42 [1518]);
assign l_41[1487]    = ( l_42 [1519]);
assign l_41[1488]    = ( l_42 [1520]);
assign l_41[1489]    = ( l_42 [1521]);
assign l_41[1490]    = ( l_42 [1522]);
assign l_41[1491]    = ( l_42 [1523]);
assign l_41[1492]    = ( l_42 [1524]);
assign l_41[1493]    = ( l_42 [1525]);
assign l_41[1494]    = ( l_42 [1526]);
assign l_41[1495]    = ( l_42 [1527]);
assign l_41[1496]    = ( l_42 [1528]);
assign l_41[1497]    = ( l_42 [1529]);
assign l_41[1498]    = ( l_42 [1530]);
assign l_41[1499]    = ( l_42 [1531]);
assign l_41[1500]    = ( l_42 [1532]);
assign l_41[1501]    = ( l_42 [1533]);
assign l_41[1502]    = ( l_42 [1534]);
assign l_41[1503]    = ( l_42 [1535]);
assign l_41[1504]    = ( l_42 [1536]);
assign l_41[1505]    = ( l_42 [1537]);
assign l_41[1506]    = ( l_42 [1538]);
assign l_41[1507]    = ( l_42 [1539]);
assign l_41[1508]    = ( l_42 [1540]);
assign l_41[1509]    = ( l_42 [1541]);
assign l_41[1510]    = ( l_42 [1542]);
assign l_41[1511]    = ( l_42 [1543]);
assign l_41[1512]    = ( l_42 [1544]);
assign l_41[1513]    = ( l_42 [1545]);
assign l_41[1514]    = ( l_42 [1546]);
assign l_41[1515]    = ( l_42 [1547]);
assign l_41[1516]    = ( l_42 [1548]);
assign l_41[1517]    = ( l_42 [1549]);
assign l_41[1518]    = ( l_42 [1550]);
assign l_41[1519]    = ( l_42 [1551]);
assign l_41[1520]    = ( l_42 [1552]);
assign l_41[1521]    = ( l_42 [1553]);
assign l_41[1522]    = ( l_42 [1554]);
assign l_41[1523]    = ( l_42 [1555]);
assign l_41[1524]    = ( l_42 [1556]);
assign l_41[1525]    = ( l_42 [1557]);
assign l_41[1526]    = ( l_42 [1558]);
assign l_41[1527]    = ( l_42 [1559]);
assign l_41[1528]    = ( l_42 [1560]);
assign l_41[1529]    = ( l_42 [1561]);
assign l_41[1530]    = ( l_42 [1562]);
assign l_41[1531]    = ( l_42 [1563]);
assign l_41[1532]    = ( l_42 [1564]);
assign l_41[1533]    = ( l_42 [1565]);
assign l_41[1534]    = ( l_42 [1566]);
assign l_41[1535]    = ( l_42 [1567]);
assign l_41[1536]    = ( l_42 [1568]);
assign l_41[1537]    = ( l_42 [1569]);
assign l_41[1538]    = ( l_42 [1570]);
assign l_41[1539]    = ( l_42 [1571]);
assign l_41[1540]    = ( l_42 [1572]);
assign l_41[1541]    = ( l_42 [1573]);
assign l_41[1542]    = ( l_42 [1574]);
assign l_41[1543]    = ( l_42 [1575]);
assign l_41[1544]    = ( l_42 [1576]);
assign l_41[1545]    = ( l_42 [1577]);
assign l_41[1546]    = ( l_42 [1578]);
assign l_41[1547]    = ( l_42 [1579]);
assign l_41[1548]    = ( l_42 [1580]);
assign l_41[1549]    = ( l_42 [1581]);
assign l_41[1550]    = ( l_42 [1582]);
assign l_41[1551]    = ( l_42 [1583]);
assign l_41[1552]    = ( l_42 [1584]);
assign l_41[1553]    = ( l_42 [1585]);
assign l_41[1554]    = ( l_42 [1586]);
assign l_41[1555]    = ( l_42 [1587]);
assign l_41[1556]    = ( l_42 [1588]);
assign l_41[1557]    = ( l_42 [1589]);
assign l_41[1558]    = ( l_42 [1590]);
assign l_41[1559]    = ( l_42 [1591]);
assign l_41[1560]    = ( l_42 [1592]);
assign l_41[1561]    = ( l_42 [1593]);
assign l_41[1562]    = ( l_42 [1594]);
assign l_41[1563]    = ( l_42 [1595]);
assign l_41[1564]    = ( l_42 [1596]);
assign l_41[1565]    = ( l_42 [1597]);
assign l_41[1566]    = ( l_42 [1598]);
assign l_41[1567]    = ( l_42 [1599]);
assign l_41[1568]    = ( l_42 [1600]);
assign l_41[1569]    = ( l_42 [1601]);
assign l_41[1570]    = ( l_42 [1602]);
assign l_41[1571]    = ( l_42 [1603]);
assign l_41[1572]    = ( l_42 [1604]);
assign l_41[1573]    = ( l_42 [1605]);
assign l_41[1574]    = ( l_42 [1606]);
assign l_41[1575]    = ( l_42 [1607]);
assign l_41[1576]    = ( l_42 [1608]);
assign l_41[1577]    = ( l_42 [1609]);
assign l_41[1578]    = ( l_42 [1610]);
assign l_41[1579]    = ( l_42 [1611]);
assign l_41[1580]    = ( l_42 [1612]);
assign l_41[1581]    = ( l_42 [1613]);
assign l_41[1582]    = ( l_42 [1614]);
assign l_41[1583]    = ( l_42 [1615]);
assign l_41[1584]    = ( l_42 [1616]);
assign l_41[1585]    = ( l_42 [1617]);
assign l_41[1586]    = ( l_42 [1618]);
assign l_41[1587]    = ( l_42 [1619]);
assign l_41[1588]    = ( l_42 [1620]);
assign l_41[1589]    = ( l_42 [1621]);
assign l_41[1590]    = ( l_42 [1622]);
assign l_41[1591]    = ( l_42 [1623]);
assign l_41[1592]    = ( l_42 [1624]);
assign l_41[1593]    = ( l_42 [1625]);
assign l_41[1594]    = ( l_42 [1626]);
assign l_41[1595]    = ( l_42 [1627]);
assign l_41[1596]    = ( l_42 [1628]);
assign l_41[1597]    = ( l_42 [1629]);
assign l_41[1598]    = ( l_42 [1630]);
assign l_41[1599]    = ( l_42 [1631]);
assign l_41[1600]    = ( l_42 [1632]);
assign l_41[1601]    = ( l_42 [1633]);
assign l_41[1602]    = ( l_42 [1634]);
assign l_41[1603]    = ( l_42 [1635]);
assign l_41[1604]    = ( l_42 [1636]);
assign l_41[1605]    = ( l_42 [1637]);
assign l_41[1606]    = ( l_42 [1638]);
assign l_41[1607]    = ( l_42 [1639]);
assign l_41[1608]    = ( l_42 [1640]);
assign l_41[1609]    = ( l_42 [1641]);
assign l_41[1610]    = ( l_42 [1642]);
assign l_41[1611]    = ( l_42 [1643]);
assign l_41[1612]    = ( l_42 [1644]);
assign l_41[1613]    = ( l_42 [1645]);
assign l_41[1614]    = ( l_42 [1646]);
assign l_41[1615]    = ( l_42 [1647]);
assign l_41[1616]    = ( l_42 [1648]);
assign l_41[1617]    = ( l_42 [1649]);
assign l_41[1618]    = ( l_42 [1650]);
assign l_41[1619]    = ( l_42 [1651]);
assign l_41[1620]    = ( l_42 [1652]);
assign l_41[1621]    = ( l_42 [1653]);
assign l_41[1622]    = ( l_42 [1654]);
assign l_41[1623]    = ( l_42 [1655]);
assign l_41[1624]    = ( l_42 [1656]);
assign l_41[1625]    = ( l_42 [1657]);
assign l_41[1626]    = ( l_42 [1658]);
assign l_41[1627]    = ( l_42 [1659]);
assign l_41[1628]    = ( l_42 [1660]);
assign l_41[1629]    = ( l_42 [1661]);
assign l_41[1630]    = ( l_42 [1662]);
assign l_41[1631]    = ( l_42 [1663]);
assign l_41[1632]    = ( l_42 [1664]);
assign l_41[1633]    = ( l_42 [1665]);
assign l_41[1634]    = ( l_42 [1666]);
assign l_41[1635]    = ( l_42 [1667]);
assign l_41[1636]    = ( l_42 [1668]);
assign l_41[1637]    = ( l_42 [1669]);
assign l_41[1638]    = ( l_42 [1670]);
assign l_41[1639]    = ( l_42 [1671]);
assign l_41[1640]    = ( l_42 [1672]);
assign l_41[1641]    = ( l_42 [1673]);
assign l_41[1642]    = ( l_42 [1674]);
assign l_41[1643]    = ( l_42 [1675]);
assign l_41[1644]    = ( l_42 [1676]);
assign l_41[1645]    = ( l_42 [1677]);
assign l_41[1646]    = ( l_42 [1678]);
assign l_41[1647]    = ( l_42 [1679]);
assign l_41[1648]    = ( l_42 [1680]);
assign l_41[1649]    = ( l_42 [1681]);
assign l_41[1650]    = ( l_42 [1682]);
assign l_41[1651]    = ( l_42 [1683]);
assign l_41[1652]    = ( l_42 [1684]);
assign l_41[1653]    = ( l_42 [1685]);
assign l_41[1654]    = ( l_42 [1686]);
assign l_41[1655]    = ( l_42 [1687]);
assign l_41[1656]    = ( l_42 [1688]);
assign l_41[1657]    = ( l_42 [1689]);
assign l_41[1658]    = ( l_42 [1690]);
assign l_41[1659]    = ( l_42 [1691]);
assign l_41[1660]    = ( l_42 [1692]);
assign l_41[1661]    = ( l_42 [1693]);
assign l_41[1662]    = ( l_42 [1694]);
assign l_41[1663]    = ( l_42 [1695]);
assign l_41[1664]    = ( l_42 [1696]);
assign l_41[1665]    = ( l_42 [1697]);
assign l_41[1666]    = ( l_42 [1698]);
assign l_41[1667]    = ( l_42 [1699]);
assign l_41[1668]    = ( l_42 [1700]);
assign l_41[1669]    = ( l_42 [1701]);
assign l_41[1670]    = ( l_42 [1702]);
assign l_41[1671]    = ( l_42 [1703]);
assign l_41[1672]    = ( l_42 [1704]);
assign l_41[1673]    = ( l_42 [1705]);
assign l_41[1674]    = ( l_42 [1706]);
assign l_41[1675]    = ( l_42 [1707]);
assign l_41[1676]    = ( l_42 [1708]);
assign l_41[1677]    = ( l_42 [1709]);
assign l_41[1678]    = ( l_42 [1710]);
assign l_41[1679]    = ( l_42 [1711]);
assign l_41[1680]    = ( l_42 [1712]);
assign l_41[1681]    = ( l_42 [1713]);
assign l_41[1682]    = ( l_42 [1714]);
assign l_41[1683]    = ( l_42 [1715]);
assign l_41[1684]    = ( l_42 [1716]);
assign l_41[1685]    = ( l_42 [1717]);
assign l_41[1686]    = ( l_42 [1718]);
assign l_41[1687]    = ( l_42 [1719]);
assign l_41[1688]    = ( l_42 [1720]);
assign l_41[1689]    = ( l_42 [1721]);
assign l_41[1690]    = ( l_42 [1722]);
assign l_41[1691]    = ( l_42 [1723]);
assign l_41[1692]    = ( l_42 [1724]);
assign l_41[1693]    = ( l_42 [1725]);
assign l_41[1694]    = ( l_42 [1726]);
assign l_41[1695]    = ( l_42 [1727]);
assign l_41[1696]    = ( l_42 [1728]);
assign l_41[1697]    = ( l_42 [1729]);
assign l_41[1698]    = ( l_42 [1730]);
assign l_41[1699]    = ( l_42 [1731]);
assign l_41[1700]    = ( l_42 [1732]);
assign l_41[1701]    = ( l_42 [1733]);
assign l_41[1702]    = ( l_42 [1734]);
assign l_41[1703]    = ( l_42 [1735]);
assign l_41[1704]    = ( l_42 [1736]);
assign l_41[1705]    = ( l_42 [1737]);
assign l_41[1706]    = ( l_42 [1738]);
assign l_41[1707]    = ( l_42 [1739]);
assign l_41[1708]    = ( l_42 [1740]);
assign l_41[1709]    = ( l_42 [1741]);
assign l_41[1710]    = ( l_42 [1742]);
assign l_41[1711]    = ( l_42 [1743]);
assign l_41[1712]    = ( l_42 [1744]);
assign l_41[1713]    = ( l_42 [1745]);
assign l_41[1714]    = ( l_42 [1746]);
assign l_41[1715]    = ( l_42 [1747]);
assign l_41[1716]    = ( l_42 [1748]);
assign l_41[1717]    = ( l_42 [1749]);
assign l_41[1718]    = ( l_42 [1750]);
assign l_41[1719]    = ( l_42 [1751]);
assign l_41[1720]    = ( l_42 [1752]);
assign l_41[1721]    = ( l_42 [1753]);
assign l_41[1722]    = ( l_42 [1754]);
assign l_41[1723]    = ( l_42 [1755]);
assign l_41[1724]    = ( l_42 [1756]);
assign l_41[1725]    = ( l_42 [1757]);
assign l_41[1726]    = ( l_42 [1758]);
assign l_41[1727]    = ( l_42 [1759]);
assign l_41[1728]    = ( l_42 [1760]);
assign l_41[1729]    = ( l_42 [1761]);
assign l_41[1730]    = ( l_42 [1762]);
assign l_41[1731]    = ( l_42 [1763]);
assign l_41[1732]    = ( l_42 [1764]);
assign l_41[1733]    = ( l_42 [1765]);
assign l_41[1734]    = ( l_42 [1766]);
assign l_41[1735]    = ( l_42 [1767]);
assign l_41[1736]    = ( l_42 [1768]);
assign l_41[1737]    = ( l_42 [1769]);
assign l_41[1738]    = ( l_42 [1770]);
assign l_41[1739]    = ( l_42 [1771]);
assign l_41[1740]    = ( l_42 [1772]);
assign l_41[1741]    = ( l_42 [1773]);
assign l_41[1742]    = ( l_42 [1774]);
assign l_41[1743]    = ( l_42 [1775]);
assign l_41[1744]    = ( l_42 [1776]);
assign l_41[1745]    = ( l_42 [1777]);
assign l_41[1746]    = ( l_42 [1778]);
assign l_41[1747]    = ( l_42 [1779]);
assign l_41[1748]    = ( l_42 [1780]);
assign l_41[1749]    = ( l_42 [1781]);
assign l_41[1750]    = ( l_42 [1782]);
assign l_41[1751]    = ( l_42 [1783]);
assign l_41[1752]    = ( l_42 [1784]);
assign l_41[1753]    = ( l_42 [1785]);
assign l_41[1754]    = ( l_42 [1786]);
assign l_41[1755]    = ( l_42 [1787]);
assign l_41[1756]    = ( l_42 [1788]);
assign l_41[1757]    = ( l_42 [1789]);
assign l_41[1758]    = ( l_42 [1790]);
assign l_41[1759]    = ( l_42 [1791]);
assign l_41[1760]    = ( l_42 [1792]);
assign l_41[1761]    = ( l_42 [1793]);
assign l_41[1762]    = ( l_42 [1794]);
assign l_41[1763]    = ( l_42 [1795]);
assign l_41[1764]    = ( l_42 [1796]);
assign l_41[1765]    = ( l_42 [1797]);
assign l_41[1766]    = ( l_42 [1798]);
assign l_41[1767]    = ( l_42 [1799]);
assign l_41[1768]    = ( l_42 [1800]);
assign l_41[1769]    = ( l_42 [1801]);
assign l_41[1770]    = ( l_42 [1802]);
assign l_41[1771]    = ( l_42 [1803]);
assign l_41[1772]    = ( l_42 [1804]);
assign l_41[1773]    = ( l_42 [1805]);
assign l_41[1774]    = ( l_42 [1806]);
assign l_41[1775]    = ( l_42 [1807]);
assign l_41[1776]    = ( l_42 [1808]);
assign l_41[1777]    = ( l_42 [1809]);
assign l_41[1778]    = ( l_42 [1810]);
assign l_41[1779]    = ( l_42 [1811]);
assign l_41[1780]    = ( l_42 [1812]);
assign l_41[1781]    = ( l_42 [1813]);
assign l_41[1782]    = ( l_42 [1814]);
assign l_41[1783]    = ( l_42 [1815]);
assign l_41[1784]    = ( l_42 [1816]);
assign l_41[1785]    = ( l_42 [1817]);
assign l_41[1786]    = ( l_42 [1818]);
assign l_41[1787]    = ( l_42 [1819]);
assign l_41[1788]    = ( l_42 [1820]);
assign l_41[1789]    = ( l_42 [1821]);
assign l_41[1790]    = ( l_42 [1822]);
assign l_41[1791]    = ( l_42 [1823]);
assign l_41[1792]    = ( l_42 [1824]);
assign l_41[1793]    = ( l_42 [1825]);
assign l_41[1794]    = ( l_42 [1826]);
assign l_41[1795]    = ( l_42 [1827]);
assign l_41[1796]    = ( l_42 [1828]);
assign l_41[1797]    = ( l_42 [1829]);
assign l_41[1798]    = ( l_42 [1830]);
assign l_41[1799]    = ( l_42 [1831]);
assign l_41[1800]    = ( l_42 [1832]);
assign l_41[1801]    = ( l_42 [1833]);
assign l_41[1802]    = ( l_42 [1834]);
assign l_41[1803]    = ( l_42 [1835]);
assign l_41[1804]    = ( l_42 [1836]);
assign l_41[1805]    = ( l_42 [1837]);
assign l_41[1806]    = ( l_42 [1838]);
assign l_41[1807]    = ( l_42 [1839]);
assign l_41[1808]    = ( l_42 [1840]);
assign l_41[1809]    = ( l_42 [1841]);
assign l_41[1810]    = ( l_42 [1842]);
assign l_41[1811]    = ( l_42 [1843]);
assign l_41[1812]    = ( l_42 [1844]);
assign l_41[1813]    = ( l_42 [1845]);
assign l_41[1814]    = ( l_42 [1846]);
assign l_41[1815]    = ( l_42 [1847]);
assign l_41[1816]    = ( l_42 [1848]);
assign l_41[1817]    = ( l_42 [1849]);
assign l_41[1818]    = ( l_42 [1850]);
assign l_41[1819]    = ( l_42 [1851]);
assign l_41[1820]    = ( l_42 [1852]);
assign l_41[1821]    = ( l_42 [1853]);
assign l_41[1822]    = ( l_42 [1854]);
assign l_41[1823]    = ( l_42 [1855]);
assign l_41[1824]    = ( l_42 [1856]);
assign l_41[1825]    = ( l_42 [1857]);
assign l_41[1826]    = ( l_42 [1858]);
assign l_41[1827]    = ( l_42 [1859]);
assign l_41[1828]    = ( l_42 [1860]);
assign l_41[1829]    = ( l_42 [1861]);
assign l_41[1830]    = ( l_42 [1862]);
assign l_41[1831]    = ( l_42 [1863]);
assign l_41[1832]    = ( l_42 [1864]);
assign l_41[1833]    = ( l_42 [1865]);
assign l_41[1834]    = ( l_42 [1866]);
assign l_41[1835]    = ( l_42 [1867]);
assign l_41[1836]    = ( l_42 [1868]);
assign l_41[1837]    = ( l_42 [1869]);
assign l_41[1838]    = ( l_42 [1870]);
assign l_41[1839]    = ( l_42 [1871]);
assign l_41[1840]    = ( l_42 [1872]);
assign l_41[1841]    = ( l_42 [1873]);
assign l_41[1842]    = ( l_42 [1874]);
assign l_41[1843]    = ( l_42 [1875]);
assign l_41[1844]    = ( l_42 [1876]);
assign l_41[1845]    = ( l_42 [1877]);
assign l_41[1846]    = ( l_42 [1878]);
assign l_41[1847]    = ( l_42 [1879]);
assign l_41[1848]    = ( l_42 [1880]);
assign l_41[1849]    = ( l_42 [1881]);
assign l_41[1850]    = ( l_42 [1882]);
assign l_41[1851]    = ( l_42 [1883]);
assign l_41[1852]    = ( l_42 [1884]);
assign l_41[1853]    = ( l_42 [1885]);
assign l_41[1854]    = ( l_42 [1886]);
assign l_41[1855]    = ( l_42 [1887]);
assign l_41[1856]    = ( l_42 [1888]);
assign l_41[1857]    = ( l_42 [1889]);
assign l_41[1858]    = ( l_42 [1890]);
assign l_41[1859]    = ( l_42 [1891]);
assign l_41[1860]    = ( l_42 [1892]);
assign l_41[1861]    = ( l_42 [1893]);
assign l_41[1862]    = ( l_42 [1894]);
assign l_41[1863]    = ( l_42 [1895]);
assign l_41[1864]    = ( l_42 [1896]);
assign l_41[1865]    = ( l_42 [1897]);
assign l_41[1866]    = ( l_42 [1898]);
assign l_41[1867]    = ( l_42 [1899]);
assign l_41[1868]    = ( l_42 [1900]);
assign l_41[1869]    = ( l_42 [1901]);
assign l_41[1870]    = ( l_42 [1902]);
assign l_41[1871]    = ( l_42 [1903]);
assign l_41[1872]    = ( l_42 [1904]);
assign l_41[1873]    = ( l_42 [1905]);
assign l_41[1874]    = ( l_42 [1906]);
assign l_41[1875]    = ( l_42 [1907]);
assign l_41[1876]    = ( l_42 [1908]);
assign l_41[1877]    = ( l_42 [1909]);
assign l_41[1878]    = ( l_42 [1910]);
assign l_41[1879]    = ( l_42 [1911]);
assign l_41[1880]    = ( l_42 [1912]);
assign l_41[1881]    = ( l_42 [1913]);
assign l_41[1882]    = ( l_42 [1914]);
assign l_41[1883]    = ( l_42 [1915]);
assign l_41[1884]    = ( l_42 [1916]);
assign l_41[1885]    = ( l_42 [1917]);
assign l_41[1886]    = ( l_42 [1918]);
assign l_41[1887]    = ( l_42 [1919]);
assign l_41[1888]    = ( l_42 [1920]);
assign l_41[1889]    = ( l_42 [1921]);
assign l_41[1890]    = ( l_42 [1922]);
assign l_41[1891]    = ( l_42 [1923]);
assign l_41[1892]    = ( l_42 [1924]);
assign l_41[1893]    = ( l_42 [1925]);
assign l_41[1894]    = ( l_42 [1926]);
assign l_41[1895]    = ( l_42 [1927]);
assign l_41[1896]    = ( l_42 [1928]);
assign l_41[1897]    = ( l_42 [1929]);
assign l_41[1898]    = ( l_42 [1930]);
assign l_41[1899]    = ( l_42 [1931]);
assign l_41[1900]    = ( l_42 [1932]);
assign l_41[1901]    = ( l_42 [1933]);
assign l_41[1902]    = ( l_42 [1934]);
assign l_41[1903]    = ( l_42 [1935]);
assign l_41[1904]    = ( l_42 [1936]);
assign l_41[1905]    = ( l_42 [1937]);
assign l_41[1906]    = ( l_42 [1938]);
assign l_41[1907]    = ( l_42 [1939]);
assign l_41[1908]    = ( l_42 [1940]);
assign l_41[1909]    = ( l_42 [1941]);
assign l_41[1910]    = ( l_42 [1942]);
assign l_41[1911]    = ( l_42 [1943]);
assign l_41[1912]    = ( l_42 [1944]);
assign l_41[1913]    = ( l_42 [1945]);
assign l_41[1914]    = ( l_42 [1946]);
assign l_41[1915]    = ( l_42 [1947]);
assign l_41[1916]    = ( l_42 [1948]);
assign l_41[1917]    = ( l_42 [1949]);
assign l_41[1918]    = ( l_42 [1950]);
assign l_41[1919]    = ( l_42 [1951]);
assign l_41[1920]    = ( l_42 [1952]);
assign l_41[1921]    = ( l_42 [1953]);
assign l_41[1922]    = ( l_42 [1954]);
assign l_41[1923]    = ( l_42 [1955]);
assign l_41[1924]    = ( l_42 [1956]);
assign l_41[1925]    = ( l_42 [1957]);
assign l_41[1926]    = ( l_42 [1958]);
assign l_41[1927]    = ( l_42 [1959]);
assign l_41[1928]    = ( l_42 [1960]);
assign l_41[1929]    = ( l_42 [1961]);
assign l_41[1930]    = ( l_42 [1962]);
assign l_41[1931]    = ( l_42 [1963]);
assign l_41[1932]    = ( l_42 [1964]);
assign l_41[1933]    = ( l_42 [1965]);
assign l_41[1934]    = ( l_42 [1966]);
assign l_41[1935]    = ( l_42 [1967]);
assign l_41[1936]    = ( l_42 [1968]);
assign l_41[1937]    = ( l_42 [1969]);
assign l_41[1938]    = ( l_42 [1970]);
assign l_41[1939]    = ( l_42 [1971]);
assign l_41[1940]    = ( l_42 [1972]);
assign l_41[1941]    = ( l_42 [1973]);
assign l_41[1942]    = ( l_42 [1974]);
assign l_41[1943]    = ( l_42 [1975]);
assign l_41[1944]    = ( l_42 [1976]);
assign l_41[1945]    = ( l_42 [1977]);
assign l_41[1946]    = ( l_42 [1978]);
assign l_41[1947]    = ( l_42 [1979]);
assign l_41[1948]    = ( l_42 [1980]);
assign l_41[1949]    = ( l_42 [1981]);
assign l_41[1950]    = ( l_42 [1982]);
assign l_41[1951]    = ( l_42 [1983]);
assign l_41[1952]    = ( l_42 [1984]);
assign l_41[1953]    = ( l_42 [1985]);
assign l_41[1954]    = ( l_42 [1986]);
assign l_41[1955]    = ( l_42 [1987]);
assign l_41[1956]    = ( l_42 [1988]);
assign l_41[1957]    = ( l_42 [1989]);
assign l_41[1958]    = ( l_42 [1990]);
assign l_41[1959]    = ( l_42 [1991]);
assign l_41[1960]    = ( l_42 [1992]);
assign l_41[1961]    = ( l_42 [1993]);
assign l_41[1962]    = ( l_42 [1994]);
assign l_41[1963]    = ( l_42 [1995]);
assign l_41[1964]    = ( l_42 [1996]);
assign l_41[1965]    = ( l_42 [1997]);
assign l_41[1966]    = ( l_42 [1998]);
assign l_41[1967]    = ( l_42 [1999]);
assign l_41[1968]    = ( l_42 [2000]);
assign l_41[1969]    = ( l_42 [2001]);
assign l_41[1970]    = ( l_42 [2002]);
assign l_41[1971]    = ( l_42 [2003]);
assign l_41[1972]    = ( l_42 [2004]);
assign l_41[1973]    = ( l_42 [2005]);
assign l_41[1974]    = ( l_42 [2006]);
assign l_41[1975]    = ( l_42 [2007]);
assign l_41[1976]    = ( l_42 [2008]);
assign l_41[1977]    = ( l_42 [2009]);
assign l_41[1978]    = ( l_42 [2010]);
assign l_41[1979]    = ( l_42 [2011]);
assign l_41[1980]    = ( l_42 [2012]);
assign l_41[1981]    = ( l_42 [2013]);
assign l_41[1982]    = ( l_42 [2014]);
assign l_41[1983]    = ( l_42 [2015]);
assign l_41[1984]    = ( l_42 [2016]);
assign l_41[1985]    = ( l_42 [2017]);
assign l_41[1986]    = ( l_42 [2018]);
assign l_41[1987]    = ( l_42 [2019]);
assign l_41[1988]    = ( l_42 [2020]);
assign l_41[1989]    = ( l_42 [2021]);
assign l_41[1990]    = ( l_42 [2022]);
assign l_41[1991]    = ( l_42 [2023]);
assign l_41[1992]    = ( l_42 [2024]);
assign l_41[1993]    = ( l_42 [2025]);
assign l_41[1994]    = ( l_42 [2026]);
assign l_41[1995]    = ( l_42 [2027]);
assign l_41[1996]    = ( l_42 [2028]);
assign l_41[1997]    = ( l_42 [2029]);
assign l_41[1998]    = ( l_42 [2030]);
assign l_41[1999]    = ( l_42 [2031]);
assign l_41[2000]    = ( l_42 [2032]);
assign l_41[2001]    = ( l_42 [2033]);
assign l_41[2002]    = ( l_42 [2034]);
assign l_41[2003]    = ( l_42 [2035]);
assign l_41[2004]    = ( l_42 [2036]);
assign l_41[2005]    = ( l_42 [2037]);
assign l_41[2006]    = ( l_42 [2038]);
assign l_41[2007]    = ( l_42 [2039]);
assign l_41[2008]    = ( l_42 [2040]);
assign l_41[2009]    = ( l_42 [2041]);
assign l_41[2010]    = ( l_42 [2042]);
assign l_41[2011]    = ( l_42 [2043]);
assign l_41[2012]    = ( l_42 [2044]);
assign l_41[2013]    = ( l_42 [2045]);
assign l_41[2014]    = ( l_42 [2046]);
assign l_41[2015]    = ( l_42 [2047]);
assign l_41[2016]    = ( l_42 [2048]);
assign l_41[2017]    = ( l_42 [2049]);
assign l_41[2018]    = ( l_42 [2050]);
assign l_41[2019]    = ( l_42 [2051]);
assign l_41[2020]    = ( l_42 [2052]);
assign l_41[2021]    = ( l_42 [2053]);
assign l_41[2022]    = ( l_42 [2054]);
assign l_41[2023]    = ( l_42 [2055]);
assign l_41[2024]    = ( l_42 [2056]);
assign l_41[2025]    = ( l_42 [2057]);
assign l_41[2026]    = ( l_42 [2058]);
assign l_41[2027]    = ( l_42 [2059]);
assign l_41[2028]    = ( l_42 [2060]);
assign l_41[2029]    = ( l_42 [2061]);
assign l_41[2030]    = ( l_42 [2062]);
assign l_41[2031]    = ( l_42 [2063]);
assign l_41[2032]    = ( l_42 [2064]);
assign l_41[2033]    = ( l_42 [2065]);
assign l_41[2034]    = ( l_42 [2066]);
assign l_41[2035]    = ( l_42 [2067]);
assign l_41[2036]    = ( l_42 [2068]);
assign l_41[2037]    = ( l_42 [2069]);
assign l_41[2038]    = ( l_42 [2070]);
assign l_41[2039]    = ( l_42 [2071]);
assign l_41[2040]    = ( l_42 [2072]);
assign l_41[2041]    = ( l_42 [2073]);
assign l_41[2042]    = ( l_42 [2074]);
assign l_41[2043]    = ( l_42 [2075]);
assign l_41[2044]    = ( l_42 [2076]);
assign l_41[2045]    = ( l_42 [2077]);
assign l_41[2046]    = ( l_42 [2078]);
assign l_41[2047]    = ( l_42 [2079]);
assign l_41[2048]    = ( l_42 [2080]);
assign l_41[2049]    = ( l_42 [2081]);
assign l_41[2050]    = ( l_42 [2082]);
assign l_41[2051]    = ( l_42 [2083]);
assign l_41[2052]    = ( l_42 [2084]);
assign l_41[2053]    = ( l_42 [2085]);
assign l_41[2054]    = ( l_42 [2086]);
assign l_41[2055]    = ( l_42 [2087]);
assign l_41[2056]    = ( l_42 [2088]);
assign l_41[2057]    = ( l_42 [2089]);
assign l_41[2058]    = ( l_42 [2090]);
assign l_41[2059]    = ( l_42 [2091]);
assign l_41[2060]    = ( l_42 [2092]);
assign l_41[2061]    = ( l_42 [2093]);
assign l_41[2062]    = ( l_42 [2094]);
assign l_41[2063]    = ( l_42 [2095]);
assign l_41[2064]    = ( l_42 [2096]);
assign l_41[2065]    = ( l_42 [2097]);
assign l_41[2066]    = ( l_42 [2098]);
assign l_41[2067]    = ( l_42 [2099]);
assign l_41[2068]    = ( l_42 [2100]);
assign l_41[2069]    = ( l_42 [2101]);
assign l_41[2070]    = ( l_42 [2102]);
assign l_41[2071]    = ( l_42 [2103]);
assign l_41[2072]    = ( l_42 [2104]);
assign l_41[2073]    = ( l_42 [2105]);
assign l_41[2074]    = ( l_42 [2106]);
assign l_41[2075]    = ( l_42 [2107]);
assign l_41[2076]    = ( l_42 [2108]);
assign l_41[2077]    = ( l_42 [2109]);
assign l_41[2078]    = ( l_42 [2110]);
assign l_41[2079]    = ( l_42 [2111]);
assign l_41[2080]    = ( l_42 [2112]);
assign l_41[2081]    = ( l_42 [2113]);
assign l_41[2082]    = ( l_42 [2114]);
assign l_41[2083]    = ( l_42 [2115]);
assign l_41[2084]    = ( l_42 [2116]);
assign l_41[2085]    = ( l_42 [2117]);
assign l_41[2086]    = ( l_42 [2118]);
assign l_41[2087]    = ( l_42 [2119]);
assign l_41[2088]    = ( l_42 [2120]);
assign l_41[2089]    = ( l_42 [2121]);
assign l_41[2090]    = ( l_42 [2122]);
assign l_41[2091]    = ( l_42 [2123]);
assign l_41[2092]    = ( l_42 [2124]);
assign l_41[2093]    = ( l_42 [2125]);
assign l_41[2094]    = ( l_42 [2126]);
assign l_41[2095]    = ( l_42 [2127]);
assign l_41[2096]    = ( l_42 [2128]);
assign l_41[2097]    = ( l_42 [2129]);
assign l_41[2098]    = ( l_42 [2130]);
assign l_41[2099]    = ( l_42 [2131]);
assign l_41[2100]    = ( l_42 [2132]);
assign l_41[2101]    = ( l_42 [2133]);
assign l_41[2102]    = ( l_42 [2134]);
assign l_41[2103]    = ( l_42 [2135]);
assign l_41[2104]    = ( l_42 [2136]);
assign l_41[2105]    = ( l_42 [2137]);
assign l_41[2106]    = ( l_42 [2138]);
assign l_41[2107]    = ( l_42 [2139]);
assign l_41[2108]    = ( l_42 [2140]);
assign l_41[2109]    = ( l_42 [2141]);
assign l_41[2110]    = ( l_42 [2142]);
assign l_41[2111]    = ( l_42 [2143]);
assign l_41[2112]    = ( l_42 [2144]);
assign l_41[2113]    = ( l_42 [2145]);
assign l_41[2114]    = ( l_42 [2146]);
assign l_41[2115]    = ( l_42 [2147]);
assign l_41[2116]    = ( l_42 [2148]);
assign l_41[2117]    = ( l_42 [2149]);
assign l_41[2118]    = ( l_42 [2150]);
assign l_41[2119]    = ( l_42 [2151]);
assign l_41[2120]    = ( l_42 [2152]);
assign l_41[2121]    = ( l_42 [2153]);
assign l_41[2122]    = ( l_42 [2154]);
assign l_41[2123]    = ( l_42 [2155]);
assign l_41[2124]    = ( l_42 [2156]);
assign l_41[2125]    = ( l_42 [2157]);
assign l_41[2126]    = ( l_42 [2158]);
assign l_41[2127]    = ( l_42 [2159]);
assign l_41[2128]    = ( l_42 [2160]);
assign l_41[2129]    = ( l_42 [2161]);
assign l_41[2130]    = ( l_42 [2162]);
assign l_41[2131]    = ( l_42 [2163]);
assign l_41[2132]    = ( l_42 [2164]);
assign l_41[2133]    = ( l_42 [2165]);
assign l_41[2134]    = ( l_42 [2166]);
assign l_41[2135]    = ( l_42 [2167]);
assign l_41[2136]    = ( l_42 [2168]);
assign l_41[2137]    = ( l_42 [2169]);
assign l_41[2138]    = ( l_42 [2170]);
assign l_41[2139]    = ( l_42 [2171]);
assign l_41[2140]    = ( l_42 [2172]);
assign l_41[2141]    = ( l_42 [2173]);
assign l_41[2142]    = ( l_42 [2174]);
assign l_41[2143]    = ( l_42 [2175]);
assign l_41[2144]    = ( l_42 [2176]);
assign l_41[2145]    = ( l_42 [2177]);
assign l_41[2146]    = ( l_42 [2178]);
assign l_41[2147]    = ( l_42 [2179]);
assign l_41[2148]    = ( l_42 [2180]);
assign l_41[2149]    = ( l_42 [2181]);
assign l_41[2150]    = ( l_42 [2182]);
assign l_41[2151]    = ( l_42 [2183]);
assign l_41[2152]    = ( l_42 [2184]);
assign l_41[2153]    = ( l_42 [2185]);
assign l_41[2154]    = ( l_42 [2186]);
assign l_41[2155]    = ( l_42 [2187]);
assign l_41[2156]    = ( l_42 [2188]);
assign l_41[2157]    = ( l_42 [2189]);
assign l_41[2158]    = ( l_42 [2190]);
assign l_41[2159]    = ( l_42 [2191]);
assign l_41[2160]    = ( l_42 [2192]);
assign l_41[2161]    = ( l_42 [2193]);
assign l_41[2162]    = ( l_42 [2194]);
assign l_41[2163]    = ( l_42 [2195]);
assign l_41[2164]    = ( l_42 [2196]);
assign l_41[2165]    = ( l_42 [2197]);
assign l_41[2166]    = ( l_42 [2198]);
assign l_41[2167]    = ( l_42 [2199]);
assign l_41[2168]    = ( l_42 [2200]);
assign l_41[2169]    = ( l_42 [2201]);
assign l_41[2170]    = ( l_42 [2202]);
assign l_41[2171]    = ( l_42 [2203]);
assign l_41[2172]    = ( l_42 [2204]);
assign l_41[2173]    = ( l_42 [2205]);
assign l_41[2174]    = ( l_42 [2206]);
assign l_41[2175]    = ( l_42 [2207]);
assign l_41[2176]    = ( l_42 [2208]);
assign l_41[2177]    = ( l_42 [2209]);
assign l_41[2178]    = ( l_42 [2210]);
assign l_41[2179]    = ( l_42 [2211]);
assign l_41[2180]    = ( l_42 [2212]);
assign l_41[2181]    = ( l_42 [2213]);
assign l_41[2182]    = ( l_42 [2214]);
assign l_41[2183]    = ( l_42 [2215]);
assign l_41[2184]    = ( l_42 [2216]);
assign l_41[2185]    = ( l_42 [2217]);
assign l_41[2186]    = ( l_42 [2218]);
assign l_41[2187]    = ( l_42 [2219]);
assign l_41[2188]    = ( l_42 [2220]);
assign l_41[2189]    = ( l_42 [2221]);
assign l_41[2190]    = ( l_42 [2222]);
assign l_41[2191]    = ( l_42 [2223]);
assign l_41[2192]    = ( l_42 [2224]);
assign l_41[2193]    = ( l_42 [2225]);
assign l_41[2194]    = ( l_42 [2226]);
assign l_41[2195]    = ( l_42 [2227]);
assign l_41[2196]    = ( l_42 [2228]);
assign l_41[2197]    = ( l_42 [2229]);
assign l_41[2198]    = ( l_42 [2230]);
assign l_41[2199]    = ( l_42 [2231]);
assign l_41[2200]    = ( l_42 [2232]);
assign l_41[2201]    = ( l_42 [2233]);
assign l_41[2202]    = ( l_42 [2234]);
assign l_41[2203]    = ( l_42 [2235]);
assign l_41[2204]    = ( l_42 [2236]);
assign l_41[2205]    = ( l_42 [2237]);
assign l_41[2206]    = ( l_42 [2238]);
assign l_41[2207]    = ( l_42 [2239]);
assign l_41[2208]    = ( l_42 [2240]);
assign l_41[2209]    = ( l_42 [2241]);
assign l_41[2210]    = ( l_42 [2242]);
assign l_41[2211]    = ( l_42 [2243]);
assign l_41[2212]    = ( l_42 [2244]);
assign l_41[2213]    = ( l_42 [2245]);
assign l_41[2214]    = ( l_42 [2246]);
assign l_41[2215]    = ( l_42 [2247]);
assign l_41[2216]    = ( l_42 [2248]);
assign l_41[2217]    = ( l_42 [2249]);
assign l_41[2218]    = ( l_42 [2250]);
assign l_41[2219]    = ( l_42 [2251]);
assign l_41[2220]    = ( l_42 [2252]);
assign l_41[2221]    = ( l_42 [2253]);
assign l_41[2222]    = ( l_42 [2254]);
assign l_41[2223]    = ( l_42 [2255]);
assign l_41[2224]    = ( l_42 [2256]);
assign l_41[2225]    = ( l_42 [2257]);
assign l_41[2226]    = ( l_42 [2258]);
assign l_41[2227]    = ( l_42 [2259]);
assign l_41[2228]    = ( l_42 [2260]);
assign l_41[2229]    = ( l_42 [2261]);
assign l_41[2230]    = ( l_42 [2262]);
assign l_41[2231]    = ( l_42 [2263]);
assign l_41[2232]    = ( l_42 [2264]);
assign l_41[2233]    = ( l_42 [2265]);
assign l_41[2234]    = ( l_42 [2266]);
assign l_41[2235]    = ( l_42 [2267]);
assign l_41[2236]    = ( l_42 [2268]);
assign l_41[2237]    = ( l_42 [2269]);
assign l_41[2238]    = ( l_42 [2270]);
assign l_41[2239]    = ( l_42 [2271]);
assign l_41[2240]    = ( l_42 [2272]);
assign l_41[2241]    = ( l_42 [2273]);
assign l_41[2242]    = ( l_42 [2274]);
assign l_41[2243]    = ( l_42 [2275]);
assign l_41[2244]    = ( l_42 [2276]);
assign l_41[2245]    = ( l_42 [2277]);
assign l_41[2246]    = ( l_42 [2278]);
assign l_41[2247]    = ( l_42 [2279]);
assign l_41[2248]    = ( l_42 [2280]);
assign l_41[2249]    = ( l_42 [2281]);
assign l_41[2250]    = ( l_42 [2282]);
assign l_41[2251]    = ( l_42 [2283]);
assign l_41[2252]    = ( l_42 [2284]);
assign l_41[2253]    = ( l_42 [2285]);
assign l_41[2254]    = ( l_42 [2286]);
assign l_41[2255]    = ( l_42 [2287]);
assign l_41[2256]    = ( l_42 [2288]);
assign l_41[2257]    = ( l_42 [2289]);
assign l_41[2258]    = ( l_42 [2290]);
assign l_41[2259]    = ( l_42 [2291]);
assign l_41[2260]    = ( l_42 [2292]);
assign l_41[2261]    = ( l_42 [2293]);
assign l_41[2262]    = ( l_42 [2294]);
assign l_41[2263]    = ( l_42 [2295]);
assign l_41[2264]    = ( l_42 [2296]);
assign l_41[2265]    = ( l_42 [2297]);
assign l_41[2266]    = ( l_42 [2298]);
assign l_41[2267]    = ( l_42 [2299]);
assign l_41[2268]    = ( l_42 [2300]);
assign l_41[2269]    = ( l_42 [2301]);
assign l_41[2270]    = ( l_42 [2302]);
assign l_41[2271]    = ( l_42 [2303]);
assign l_41[2272]    = ( l_42 [2304]);
assign l_41[2273]    = ( l_42 [2305]);
assign l_41[2274]    = ( l_42 [2306]);
assign l_41[2275]    = ( l_42 [2307]);
assign l_41[2276]    = ( l_42 [2308]);
assign l_41[2277]    = ( l_42 [2309]);
assign l_41[2278]    = ( l_42 [2310]);
assign l_41[2279]    = ( l_42 [2311]);
assign l_41[2280]    = ( l_42 [2312]);
assign l_41[2281]    = ( l_42 [2313]);
assign l_41[2282]    = ( l_42 [2314]);
assign l_41[2283]    = ( l_42 [2315]);
assign l_41[2284]    = ( l_42 [2316]);
assign l_41[2285]    = ( l_42 [2317]);
assign l_41[2286]    = ( l_42 [2318]);
assign l_41[2287]    = ( l_42 [2319]);
assign l_41[2288]    = ( l_42 [2320]);
assign l_41[2289]    = ( l_42 [2321]);
assign l_41[2290]    = ( l_42 [2322]);
assign l_41[2291]    = ( l_42 [2323]);
assign l_41[2292]    = ( l_42 [2324]);
assign l_41[2293]    = ( l_42 [2325]);
assign l_41[2294]    = ( l_42 [2326]);
assign l_41[2295]    = ( l_42 [2327]);
assign l_41[2296]    = ( l_42 [2328]);
assign l_41[2297]    = ( l_42 [2329]);
assign l_41[2298]    = ( l_42 [2330]);
assign l_41[2299]    = ( l_42 [2331]);
assign l_41[2300]    = ( l_42 [2332]);
assign l_41[2301]    = ( l_42 [2333]);
assign l_41[2302]    = ( l_42 [2334]);
assign l_41[2303]    = ( l_42 [2335]);
assign l_41[2304]    = ( l_42 [2336]);
assign l_41[2305]    = ( l_42 [2337]);
assign l_41[2306]    = ( l_42 [2338]);
assign l_41[2307]    = ( l_42 [2339]);
assign l_41[2308]    = ( l_42 [2340]);
assign l_41[2309]    = ( l_42 [2341]);
assign l_41[2310]    = ( l_42 [2342]);
assign l_41[2311]    = ( l_42 [2343]);
assign l_41[2312]    = ( l_42 [2344]);
assign l_41[2313]    = ( l_42 [2345]);
assign l_41[2314]    = ( l_42 [2346]);
assign l_41[2315]    = ( l_42 [2347]);
assign l_41[2316]    = ( l_42 [2348]);
assign l_41[2317]    = ( l_42 [2349]);
assign l_41[2318]    = ( l_42 [2350]);
assign l_41[2319]    = ( l_42 [2351]);
assign l_41[2320]    = ( l_42 [2352]);
assign l_41[2321]    = ( l_42 [2353]);
assign l_41[2322]    = ( l_42 [2354]);
assign l_41[2323]    = ( l_42 [2355]);
assign l_41[2324]    = ( l_42 [2356]);
assign l_41[2325]    = ( l_42 [2357]);
assign l_41[2326]    = ( l_42 [2358]);
assign l_41[2327]    = ( l_42 [2359]);
assign l_41[2328]    = ( l_42 [2360]);
assign l_41[2329]    = ( l_42 [2361]);
assign l_41[2330]    = ( l_42 [2362]);
assign l_41[2331]    = ( l_42 [2363]);
assign l_41[2332]    = ( l_42 [2364]);
assign l_41[2333]    = ( l_42 [2365]);
assign l_41[2334]    = ( l_42 [2366]);
assign l_41[2335]    = ( l_42 [2367]);
assign l_41[2336]    = ( l_42 [2368]);
assign l_41[2337]    = ( l_42 [2369]);
assign l_41[2338]    = ( l_42 [2370]);
assign l_41[2339]    = ( l_42 [2371]);
assign l_41[2340]    = ( l_42 [2372]);
assign l_41[2341]    = ( l_42 [2373]);
assign l_41[2342]    = ( l_42 [2374]);
assign l_41[2343]    = ( l_42 [2375]);
assign l_41[2344]    = ( l_42 [2376]);
assign l_41[2345]    = ( l_42 [2377]);
assign l_41[2346]    = ( l_42 [2378]);
assign l_41[2347]    = ( l_42 [2379]);
assign l_41[2348]    = ( l_42 [2380]);
assign l_41[2349]    = ( l_42 [2381]);
assign l_41[2350]    = ( l_42 [2382]);
assign l_41[2351]    = ( l_42 [2383]);
assign l_41[2352]    = ( l_42 [2384]);
assign l_41[2353]    = ( l_42 [2385]);
assign l_41[2354]    = ( l_42 [2386]);
assign l_41[2355]    = ( l_42 [2387]);
assign l_41[2356]    = ( l_42 [2388]);
assign l_41[2357]    = ( l_42 [2389]);
assign l_41[2358]    = ( l_42 [2390]);
assign l_41[2359]    = ( l_42 [2391]);
assign l_41[2360]    = ( l_42 [2392]);
assign l_41[2361]    = ( l_42 [2393]);
assign l_41[2362]    = ( l_42 [2394]);
assign l_41[2363]    = ( l_42 [2395]);
assign l_41[2364]    = ( l_42 [2396]);
assign l_41[2365]    = ( l_42 [2397]);
assign l_41[2366]    = ( l_42 [2398]);
assign l_41[2367]    = ( l_42 [2399]);
assign l_41[2368]    = ( l_42 [2400]);
assign l_41[2369]    = ( l_42 [2401]);
assign l_41[2370]    = ( l_42 [2402]);
assign l_41[2371]    = ( l_42 [2403]);
assign l_41[2372]    = ( l_42 [2404]);
assign l_41[2373]    = ( l_42 [2405]);
assign l_41[2374]    = ( l_42 [2406]);
assign l_41[2375]    = ( l_42 [2407]);
assign l_41[2376]    = ( l_42 [2408]);
assign l_41[2377]    = ( l_42 [2409]);
assign l_41[2378]    = ( l_42 [2410]);
assign l_41[2379]    = ( l_42 [2411]);
assign l_41[2380]    = ( l_42 [2412]);
assign l_41[2381]    = ( l_42 [2413]);
assign l_41[2382]    = ( l_42 [2414]);
assign l_41[2383]    = ( l_42 [2415]);
assign l_41[2384]    = ( l_42 [2416]);
assign l_41[2385]    = ( l_42 [2417]);
assign l_41[2386]    = ( l_42 [2418]);
assign l_41[2387]    = ( l_42 [2419]);
assign l_41[2388]    = ( l_42 [2420]);
assign l_41[2389]    = ( l_42 [2421]);
assign l_41[2390]    = ( l_42 [2422]);
assign l_41[2391]    = ( l_42 [2423]);
assign l_41[2392]    = ( l_42 [2424]);
assign l_41[2393]    = ( l_42 [2425]);
assign l_41[2394]    = ( l_42 [2426]);
assign l_41[2395]    = ( l_42 [2427]);
assign l_41[2396]    = ( l_42 [2428]);
assign l_41[2397]    = ( l_42 [2429]);
assign l_41[2398]    = ( l_42 [2430]);
assign l_41[2399]    = ( l_42 [2431]);
assign l_41[2400]    = ( l_42 [2432]);
assign l_41[2401]    = ( l_42 [2433]);
assign l_41[2402]    = ( l_42 [2434]);
assign l_41[2403]    = ( l_42 [2435]);
assign l_41[2404]    = ( l_42 [2436]);
assign l_41[2405]    = ( l_42 [2437]);
assign l_41[2406]    = ( l_42 [2438]);
assign l_41[2407]    = ( l_42 [2439]);
assign l_41[2408]    = ( l_42 [2440]);
assign l_41[2409]    = ( l_42 [2441]);
assign l_41[2410]    = ( l_42 [2442]);
assign l_41[2411]    = ( l_42 [2443]);
assign l_41[2412]    = ( l_42 [2444]);
assign l_41[2413]    = ( l_42 [2445]);
assign l_41[2414]    = ( l_42 [2446]);
assign l_41[2415]    = ( l_42 [2447]);
assign l_41[2416]    = ( l_42 [2448]);
assign l_41[2417]    = ( l_42 [2449]);
assign l_41[2418]    = ( l_42 [2450]);
assign l_41[2419]    = ( l_42 [2451]);
assign l_41[2420]    = ( l_42 [2452]);
assign l_41[2421]    = ( l_42 [2453]);
assign l_41[2422]    = ( l_42 [2454]);
assign l_41[2423]    = ( l_42 [2455]);
assign l_41[2424]    = ( l_42 [2456]);
assign l_41[2425]    = ( l_42 [2457]);
assign l_41[2426]    = ( l_42 [2458]);
assign l_41[2427]    = ( l_42 [2459]);
assign l_41[2428]    = ( l_42 [2460]);
assign l_41[2429]    = ( l_42 [2461]);
assign l_41[2430]    = ( l_42 [2462]);
assign l_41[2431]    = ( l_42 [2463]);
assign l_41[2432]    = ( l_42 [2464]);
assign l_41[2433]    = ( l_42 [2465]);
assign l_41[2434]    = ( l_42 [2466]);
assign l_41[2435]    = ( l_42 [2467]);
assign l_41[2436]    = ( l_42 [2468]);
assign l_41[2437]    = ( l_42 [2469]);
assign l_41[2438]    = ( l_42 [2470]);
assign l_41[2439]    = ( l_42 [2471]);
assign l_41[2440]    = ( l_42 [2472]);
assign l_41[2441]    = ( l_42 [2473]);
assign l_41[2442]    = ( l_42 [2474]);
assign l_41[2443]    = ( l_42 [2475]);
assign l_41[2444]    = ( l_42 [2476]);
assign l_41[2445]    = ( l_42 [2477]);
assign l_41[2446]    = ( l_42 [2478]);
assign l_41[2447]    = ( l_42 [2479]);
assign l_41[2448]    = ( l_42 [2480]);
assign l_41[2449]    = ( l_42 [2481]);
assign l_41[2450]    = ( l_42 [2482]);
assign l_41[2451]    = ( l_42 [2483]);
assign l_41[2452]    = ( l_42 [2484]);
assign l_41[2453]    = ( l_42 [2485]);
assign l_41[2454]    = ( l_42 [2486]);
assign l_41[2455]    = ( l_42 [2487]);
assign l_41[2456]    = ( l_42 [2488]);
assign l_41[2457]    = ( l_42 [2489]);
assign l_41[2458]    = ( l_42 [2490]);
assign l_41[2459]    = ( l_42 [2491]);
assign l_41[2460]    = ( l_42 [2492]);
assign l_41[2461]    = ( l_42 [2493]);
assign l_41[2462]    = ( l_42 [2494]);
assign l_41[2463]    = ( l_42 [2495]);
assign l_41[2464]    = ( l_42 [2496]);
assign l_41[2465]    = ( l_42 [2497]);
assign l_41[2466]    = ( l_42 [2498]);
assign l_41[2467]    = ( l_42 [2499]);
assign l_41[2468]    = ( l_42 [2500]);
assign l_41[2469]    = ( l_42 [2501]);
assign l_41[2470]    = ( l_42 [2502]);
assign l_41[2471]    = ( l_42 [2503]);
assign l_41[2472]    = ( l_42 [2504]);
assign l_41[2473]    = ( l_42 [2505]);
assign l_41[2474]    = ( l_42 [2506]);
assign l_41[2475]    = ( l_42 [2507]);
assign l_41[2476]    = ( l_42 [2508]);
assign l_41[2477]    = ( l_42 [2509]);
assign l_41[2478]    = ( l_42 [2510]);
assign l_41[2479]    = ( l_42 [2511]);
assign l_41[2480]    = ( l_42 [2512]);
assign l_41[2481]    = ( l_42 [2513]);
assign l_41[2482]    = ( l_42 [2514]);
assign l_41[2483]    = ( l_42 [2515]);
assign l_41[2484]    = ( l_42 [2516]);
assign l_41[2485]    = ( l_42 [2517]);
assign l_41[2486]    = ( l_42 [2518]);
assign l_41[2487]    = ( l_42 [2519]);
assign l_41[2488]    = ( l_42 [2520]);
assign l_41[2489]    = ( l_42 [2521]);
assign l_41[2490]    = ( l_42 [2522]);
assign l_41[2491]    = ( l_42 [2523]);
assign l_41[2492]    = ( l_42 [2524]);
assign l_41[2493]    = ( l_42 [2525]);
assign l_41[2494]    = ( l_42 [2526]);
assign l_41[2495]    = ( l_42 [2527]);
assign l_41[2496]    = ( l_42 [2528]);
assign l_41[2497]    = ( l_42 [2529]);
assign l_41[2498]    = ( l_42 [2530]);
assign l_41[2499]    = ( l_42 [2531]);
assign l_41[2500]    = ( l_42 [2532]);
assign l_41[2501]    = ( l_42 [2533]);
assign l_41[2502]    = ( l_42 [2534]);
assign l_41[2503]    = ( l_42 [2535]);
assign l_41[2504]    = ( l_42 [2536]);
assign l_41[2505]    = ( l_42 [2537]);
assign l_41[2506]    = ( l_42 [2538]);
assign l_41[2507]    = ( l_42 [2539]);
assign l_41[2508]    = ( l_42 [2540]);
assign l_41[2509]    = ( l_42 [2541]);
assign l_41[2510]    = ( l_42 [2542]);
assign l_41[2511]    = ( l_42 [2543]);
assign l_41[2512]    = ( l_42 [2544]);
assign l_41[2513]    = ( l_42 [2545]);
assign l_41[2514]    = ( l_42 [2546]);
assign l_41[2515]    = ( l_42 [2547]);
assign l_41[2516]    = ( l_42 [2548]);
assign l_41[2517]    = ( l_42 [2549]);
assign l_41[2518]    = ( l_42 [2550]);
assign l_41[2519]    = ( l_42 [2551]);
assign l_41[2520]    = ( l_42 [2552]);
assign l_41[2521]    = ( l_42 [2553]);
assign l_41[2522]    = ( l_42 [2554]);
assign l_41[2523]    = ( l_42 [2555]);
assign l_41[2524]    = ( l_42 [2556]);
assign l_41[2525]    = ( l_42 [2557]);
assign l_41[2526]    = ( l_42 [2558]);
assign l_41[2527]    = ( l_42 [2559]);
assign l_41[2528]    = ( l_42 [2560]);
assign l_41[2529]    = ( l_42 [2561]);
assign l_41[2530]    = ( l_42 [2562]);
assign l_41[2531]    = ( l_42 [2563]);
assign l_41[2532]    = ( l_42 [2564]);
assign l_41[2533]    = ( l_42 [2565]);
assign l_41[2534]    = ( l_42 [2566]);
assign l_41[2535]    = ( l_42 [2567]);
assign l_41[2536]    = ( l_42 [2568]);
assign l_41[2537]    = ( l_42 [2569]);
assign l_41[2538]    = ( l_42 [2570]);
assign l_41[2539]    = ( l_42 [2571]);
assign l_41[2540]    = ( l_42 [2572]);
assign l_41[2541]    = ( l_42 [2573]);
assign l_41[2542]    = ( l_42 [2574]);
assign l_41[2543]    = ( l_42 [2575]);
assign l_41[2544]    = ( l_42 [2576]);
assign l_41[2545]    = ( l_42 [2577]);
assign l_41[2546]    = ( l_42 [2578]);
assign l_41[2547]    = ( l_42 [2579]);
assign l_41[2548]    = ( l_42 [2580]);
assign l_41[2549]    = ( l_42 [2581]);
assign l_41[2550]    = ( l_42 [2582]);
assign l_41[2551]    = ( l_42 [2583]);
assign l_41[2552]    = ( l_42 [2584]);
assign l_41[2553]    = ( l_42 [2585]);
assign l_41[2554]    = ( l_42 [2586]);
assign l_41[2555]    = ( l_42 [2587]);
assign l_41[2556]    = ( l_42 [2588]);
assign l_41[2557]    = ( l_42 [2589]);
assign l_41[2558]    = ( l_42 [2590]);
assign l_41[2559]    = ( l_42 [2591]);
assign l_41[2560]    = ( l_42 [2592]);
assign l_41[2561]    = ( l_42 [2593]);
assign l_41[2562]    = ( l_42 [2594]);
assign l_41[2563]    = ( l_42 [2595]);
assign l_41[2564]    = ( l_42 [2596]);
assign l_41[2565]    = ( l_42 [2597]);
assign l_41[2566]    = ( l_42 [2598]);
assign l_41[2567]    = ( l_42 [2599]);
assign l_41[2568]    = ( l_42 [2600]);
assign l_41[2569]    = ( l_42 [2601]);
assign l_41[2570]    = ( l_42 [2602]);
assign l_41[2571]    = ( l_42 [2603]);
assign l_41[2572]    = ( l_42 [2604]);
assign l_41[2573]    = ( l_42 [2605]);
assign l_41[2574]    = ( l_42 [2606]);
assign l_41[2575]    = ( l_42 [2607]);
assign l_41[2576]    = ( l_42 [2608]);
assign l_41[2577]    = ( l_42 [2609]);
assign l_41[2578]    = ( l_42 [2610]);
assign l_41[2579]    = ( l_42 [2611]);
assign l_41[2580]    = ( l_42 [2612]);
assign l_41[2581]    = ( l_42 [2613]);
assign l_41[2582]    = ( l_42 [2614]);
assign l_41[2583]    = ( l_42 [2615]);
assign l_41[2584]    = ( l_42 [2616]);
assign l_41[2585]    = ( l_42 [2617]);
assign l_41[2586]    = ( l_42 [2618]);
assign l_41[2587]    = ( l_42 [2619]);
assign l_41[2588]    = ( l_42 [2620]);
assign l_41[2589]    = ( l_42 [2621]);
assign l_41[2590]    = ( l_42 [2622]);
assign l_41[2591]    = ( l_42 [2623]);
assign l_41[2592]    = ( l_42 [2624]);
assign l_41[2593]    = ( l_42 [2625]);
assign l_41[2594]    = ( l_42 [2626]);
assign l_41[2595]    = ( l_42 [2627]);
assign l_41[2596]    = ( l_42 [2628]);
assign l_41[2597]    = ( l_42 [2629]);
assign l_41[2598]    = ( l_42 [2630]);
assign l_41[2599]    = ( l_42 [2631]);
assign l_41[2600]    = ( l_42 [2632]);
assign l_41[2601]    = ( l_42 [2633]);
assign l_41[2602]    = ( l_42 [2634]);
assign l_41[2603]    = ( l_42 [2635]);
assign l_41[2604]    = ( l_42 [2636]);
assign l_41[2605]    = ( l_42 [2637]);
assign l_41[2606]    = ( l_42 [2638]);
assign l_41[2607]    = ( l_42 [2639]);
assign l_41[2608]    = ( l_42 [2640]);
assign l_41[2609]    = ( l_42 [2641]);
assign l_41[2610]    = ( l_42 [2642]);
assign l_41[2611]    = ( l_42 [2643]);
assign l_41[2612]    = ( l_42 [2644]);
assign l_41[2613]    = ( l_42 [2645]);
assign l_41[2614]    = ( l_42 [2646]);
assign l_41[2615]    = ( l_42 [2647]);
assign l_41[2616]    = ( l_42 [2648]);
assign l_41[2617]    = ( l_42 [2649]);
assign l_41[2618]    = ( l_42 [2650]);
assign l_41[2619]    = ( l_42 [2651]);
assign l_41[2620]    = ( l_42 [2652]);
assign l_41[2621]    = ( l_42 [2653]);
assign l_41[2622]    = ( l_42 [2654]);
assign l_41[2623]    = ( l_42 [2655]);
assign l_41[2624]    = ( l_42 [2656]);
assign l_41[2625]    = ( l_42 [2657]);
assign l_41[2626]    = ( l_42 [2658]);
assign l_41[2627]    = ( l_42 [2659]);
assign l_41[2628]    = ( l_42 [2660]);
assign l_41[2629]    = ( l_42 [2661]);
assign l_41[2630]    = ( l_42 [2662]);
assign l_41[2631]    = ( l_42 [2663]);
assign l_41[2632]    = ( l_42 [2664]);
assign l_41[2633]    = ( l_42 [2665]);
assign l_41[2634]    = ( l_42 [2666]);
assign l_41[2635]    = ( l_42 [2667]);
assign l_41[2636]    = ( l_42 [2668]);
assign l_41[2637]    = ( l_42 [2669]);
assign l_41[2638]    = ( l_42 [2670]);
assign l_41[2639]    = ( l_42 [2671]);
assign l_41[2640]    = ( l_42 [2672]);
assign l_41[2641]    = ( l_42 [2673]);
assign l_41[2642]    = ( l_42 [2674]);
assign l_41[2643]    = ( l_42 [2675]);
assign l_41[2644]    = ( l_42 [2676]);
assign l_41[2645]    = ( l_42 [2677]);
assign l_41[2646]    = ( l_42 [2678]);
assign l_41[2647]    = ( l_42 [2679]);
assign l_41[2648]    = ( l_42 [2680]);
assign l_41[2649]    = ( l_42 [2681]);
assign l_41[2650]    = ( l_42 [2682]);
assign l_41[2651]    = ( l_42 [2683]);
assign l_41[2652]    = ( l_42 [2684]);
assign l_41[2653]    = ( l_42 [2685]);
assign l_41[2654]    = ( l_42 [2686]);
assign l_41[2655]    = ( l_42 [2687]);
assign l_41[2656]    = ( l_42 [2688]);
assign l_41[2657]    = ( l_42 [2689]);
assign l_41[2658]    = ( l_42 [2690]);
assign l_41[2659]    = ( l_42 [2691]);
assign l_41[2660]    = ( l_42 [2692]);
assign l_41[2661]    = ( l_42 [2693]);
assign l_41[2662]    = ( l_42 [2694]);
assign l_41[2663]    = ( l_42 [2695]);
assign l_41[2664]    = ( l_42 [2696]);
assign l_41[2665]    = ( l_42 [2697]);
assign l_41[2666]    = ( l_42 [2698]);
assign l_41[2667]    = ( l_42 [2699]);
assign l_41[2668]    = ( l_42 [2700]);
assign l_41[2669]    = ( l_42 [2701]);
assign l_41[2670]    = ( l_42 [2702]);
assign l_41[2671]    = ( l_42 [2703]);
assign l_41[2672]    = ( l_42 [2704]);
assign l_41[2673]    = ( l_42 [2705]);
assign l_41[2674]    = ( l_42 [2706]);
assign l_41[2675]    = ( l_42 [2707]);
assign l_41[2676]    = ( l_42 [2708]);
assign l_41[2677]    = ( l_42 [2709]);
assign l_41[2678]    = ( l_42 [2710]);
assign l_41[2679]    = ( l_42 [2711]);
assign l_41[2680]    = ( l_42 [2712]);
assign l_41[2681]    = ( l_42 [2713]);
assign l_41[2682]    = ( l_42 [2714]);
assign l_41[2683]    = ( l_42 [2715]);
assign l_41[2684]    = ( l_42 [2716]);
assign l_41[2685]    = ( l_42 [2717]);
assign l_41[2686]    = ( l_42 [2718]);
assign l_41[2687]    = ( l_42 [2719]);
assign l_41[2688]    = ( l_42 [2720]);
assign l_41[2689]    = ( l_42 [2721]);
assign l_41[2690]    = ( l_42 [2722]);
assign l_41[2691]    = ( l_42 [2723]);
assign l_41[2692]    = ( l_42 [2724]);
assign l_41[2693]    = ( l_42 [2725]);
assign l_41[2694]    = ( l_42 [2726]);
assign l_41[2695]    = ( l_42 [2727]);
assign l_41[2696]    = ( l_42 [2728]);
assign l_41[2697]    = ( l_42 [2729]);
assign l_41[2698]    = ( l_42 [2730]);
assign l_41[2699]    = ( l_42 [2731]);
assign l_41[2700]    = ( l_42 [2732]);
assign l_41[2701]    = ( l_42 [2733]);
assign l_41[2702]    = ( l_42 [2734]);
assign l_41[2703]    = ( l_42 [2735]);
assign l_41[2704]    = ( l_42 [2736]);
assign l_41[2705]    = ( l_42 [2737]);
assign l_41[2706]    = ( l_42 [2738]);
assign l_41[2707]    = ( l_42 [2739]);
assign l_41[2708]    = ( l_42 [2740]);
assign l_41[2709]    = ( l_42 [2741]);
assign l_41[2710]    = ( l_42 [2742]);
assign l_41[2711]    = ( l_42 [2743]);
assign l_41[2712]    = ( l_42 [2744]);
assign l_41[2713]    = ( l_42 [2745]);
assign l_41[2714]    = ( l_42 [2746]);
assign l_41[2715]    = ( l_42 [2747]);
assign l_41[2716]    = ( l_42 [2748]);
assign l_41[2717]    = ( l_42 [2749]);
assign l_41[2718]    = ( l_42 [2750]);
assign l_41[2719]    = ( l_42 [2751]);
assign l_41[2720]    = ( l_42 [2752]);
assign l_41[2721]    = ( l_42 [2753]);
assign l_41[2722]    = ( l_42 [2754]);
assign l_41[2723]    = ( l_42 [2755]);
assign l_41[2724]    = ( l_42 [2756]);
assign l_41[2725]    = ( l_42 [2757]);
assign l_41[2726]    = ( l_42 [2758]);
assign l_41[2727]    = ( l_42 [2759]);
assign l_41[2728]    = ( l_42 [2760]);
assign l_41[2729]    = ( l_42 [2761]);
assign l_41[2730]    = ( l_42 [2762]);
assign l_41[2731]    = ( l_42 [2763]);
assign l_41[2732]    = ( l_42 [2764]);
assign l_41[2733]    = ( l_42 [2765]);
assign l_41[2734]    = ( l_42 [2766]);
assign l_41[2735]    = ( l_42 [2767]);
assign l_41[2736]    = ( l_42 [2768]);
assign l_41[2737]    = ( l_42 [2769]);
assign l_41[2738]    = ( l_42 [2770]);
assign l_41[2739]    = ( l_42 [2771]);
assign l_41[2740]    = ( l_42 [2772]);
assign l_41[2741]    = ( l_42 [2773]);
assign l_41[2742]    = ( l_42 [2774]);
assign l_41[2743]    = ( l_42 [2775]);
assign l_41[2744]    = ( l_42 [2776]);
assign l_41[2745]    = ( l_42 [2777]);
assign l_41[2746]    = ( l_42 [2778]);
assign l_41[2747]    = ( l_42 [2779]);
assign l_41[2748]    = ( l_42 [2780]);
assign l_41[2749]    = ( l_42 [2781]);
assign l_41[2750]    = ( l_42 [2782]);
assign l_41[2751]    = ( l_42 [2783]);
assign l_41[2752]    = ( l_42 [2784]);
assign l_41[2753]    = ( l_42 [2785]);
assign l_41[2754]    = ( l_42 [2786]);
assign l_41[2755]    = ( l_42 [2787]);
assign l_41[2756]    = ( l_42 [2788]);
assign l_41[2757]    = ( l_42 [2789]);
assign l_41[2758]    = ( l_42 [2790]);
assign l_41[2759]    = ( l_42 [2791]);
assign l_41[2760]    = ( l_42 [2792]);
assign l_41[2761]    = ( l_42 [2793]);
assign l_41[2762]    = ( l_42 [2794]);
assign l_41[2763]    = ( l_42 [2795]);
assign l_41[2764]    = ( l_42 [2796]);
assign l_41[2765]    = ( l_42 [2797]);
assign l_41[2766]    = ( l_42 [2798]);
assign l_41[2767]    = ( l_42 [2799]);
assign l_41[2768]    = ( l_42 [2800]);
assign l_41[2769]    = ( l_42 [2801]);
assign l_41[2770]    = ( l_42 [2802]);
assign l_41[2771]    = ( l_42 [2803]);
assign l_41[2772]    = ( l_42 [2804]);
assign l_41[2773]    = ( l_42 [2805]);
assign l_41[2774]    = ( l_42 [2806]);
assign l_41[2775]    = ( l_42 [2807]);
assign l_41[2776]    = ( l_42 [2808]);
assign l_41[2777]    = ( l_42 [2809]);
assign l_41[2778]    = ( l_42 [2810]);
assign l_41[2779]    = ( l_42 [2811]);
assign l_41[2780]    = ( l_42 [2812]);
assign l_41[2781]    = ( l_42 [2813]);
assign l_41[2782]    = ( l_42 [2814]);
assign l_41[2783]    = ( l_42 [2815]);
assign l_41[2784]    = ( l_42 [2816]);
assign l_41[2785]    = ( l_42 [2817]);
assign l_41[2786]    = ( l_42 [2818]);
assign l_41[2787]    = ( l_42 [2819]);
assign l_41[2788]    = ( l_42 [2820]);
assign l_41[2789]    = ( l_42 [2821]);
assign l_41[2790]    = ( l_42 [2822]);
assign l_41[2791]    = ( l_42 [2823]);
assign l_41[2792]    = ( l_42 [2824]);
assign l_41[2793]    = ( l_42 [2825]);
assign l_41[2794]    = ( l_42 [2826]);
assign l_41[2795]    = ( l_42 [2827]);
assign l_41[2796]    = ( l_42 [2828]);
assign l_41[2797]    = ( l_42 [2829]);
assign l_41[2798]    = ( l_42 [2830]);
assign l_41[2799]    = ( l_42 [2831]);
assign l_41[2800]    = ( l_42 [2832]);
assign l_41[2801]    = ( l_42 [2833]);
assign l_41[2802]    = ( l_42 [2834]);
assign l_41[2803]    = ( l_42 [2835]);
assign l_41[2804]    = ( l_42 [2836]);
assign l_41[2805]    = ( l_42 [2837]);
assign l_41[2806]    = ( l_42 [2838]);
assign l_41[2807]    = ( l_42 [2839]);
assign l_41[2808]    = ( l_42 [2840]);
assign l_41[2809]    = ( l_42 [2841]);
assign l_41[2810]    = ( l_42 [2842]);
assign l_41[2811]    = ( l_42 [2843]);
assign l_41[2812]    = ( l_42 [2844]);
assign l_41[2813]    = ( l_42 [2845]);
assign l_41[2814]    = ( l_42 [2846]);
assign l_41[2815]    = ( l_42 [2847]);
assign l_41[2816]    = ( l_42 [2848]);
assign l_41[2817]    = ( l_42 [2849]);
assign l_41[2818]    = ( l_42 [2850]);
assign l_41[2819]    = ( l_42 [2851]);
assign l_41[2820]    = ( l_42 [2852]);
assign l_41[2821]    = ( l_42 [2853]);
assign l_41[2822]    = ( l_42 [2854]);
assign l_41[2823]    = ( l_42 [2855]);
assign l_41[2824]    = ( l_42 [2856]);
assign l_41[2825]    = ( l_42 [2857]);
assign l_41[2826]    = ( l_42 [2858]);
assign l_41[2827]    = ( l_42 [2859]);
assign l_41[2828]    = ( l_42 [2860]);
assign l_41[2829]    = ( l_42 [2861]);
assign l_41[2830]    = ( l_42 [2862]);
assign l_41[2831]    = ( l_42 [2863]);
assign l_41[2832]    = ( l_42 [2864]);
assign l_41[2833]    = ( l_42 [2865]);
assign l_41[2834]    = ( l_42 [2866]);
assign l_41[2835]    = ( l_42 [2867]);
assign l_41[2836]    = ( l_42 [2868]);
assign l_41[2837]    = ( l_42 [2869]);
assign l_41[2838]    = ( l_42 [2870]);
assign l_41[2839]    = ( l_42 [2871]);
assign l_41[2840]    = ( l_42 [2872]);
assign l_41[2841]    = ( l_42 [2873]);
assign l_41[2842]    = ( l_42 [2874]);
assign l_41[2843]    = ( l_42 [2875]);
assign l_41[2844]    = ( l_42 [2876]);
assign l_41[2845]    = ( l_42 [2877]);
assign l_41[2846]    = ( l_42 [2878]);
assign l_41[2847]    = ( l_42 [2879]);
assign l_41[2848]    = ( l_42 [2880]);
assign l_41[2849]    = ( l_42 [2881]);
assign l_41[2850]    = ( l_42 [2882]);
assign l_41[2851]    = ( l_42 [2883]);
assign l_41[2852]    = ( l_42 [2884]);
assign l_41[2853]    = ( l_42 [2885]);
assign l_41[2854]    = ( l_42 [2886]);
assign l_41[2855]    = ( l_42 [2887]);
assign l_41[2856]    = ( l_42 [2888]);
assign l_41[2857]    = ( l_42 [2889]);
assign l_41[2858]    = ( l_42 [2890]);
assign l_41[2859]    = ( l_42 [2891]);
assign l_41[2860]    = ( l_42 [2892]);
assign l_41[2861]    = ( l_42 [2893]);
assign l_41[2862]    = ( l_42 [2894]);
assign l_41[2863]    = ( l_42 [2895]);
assign l_41[2864]    = ( l_42 [2896]);
assign l_41[2865]    = ( l_42 [2897]);
assign l_41[2866]    = ( l_42 [2898]);
assign l_41[2867]    = ( l_42 [2899]);
assign l_41[2868]    = ( l_42 [2900]);
assign l_41[2869]    = ( l_42 [2901]);
assign l_41[2870]    = ( l_42 [2902]);
assign l_41[2871]    = ( l_42 [2903]);
assign l_41[2872]    = ( l_42 [2904]);
assign l_41[2873]    = ( l_42 [2905]);
assign l_41[2874]    = ( l_42 [2906]);
assign l_41[2875]    = ( l_42 [2907]);
assign l_41[2876]    = ( l_42 [2908]);
assign l_41[2877]    = ( l_42 [2909]);
assign l_41[2878]    = ( l_42 [2910]);
assign l_41[2879]    = ( l_42 [2911]);
assign l_41[2880]    = ( l_42 [2912]);
assign l_41[2881]    = ( l_42 [2913]);
assign l_41[2882]    = ( l_42 [2914]);
assign l_41[2883]    = ( l_42 [2915]);
assign l_41[2884]    = ( l_42 [2916]);
assign l_41[2885]    = ( l_42 [2917]);
assign l_41[2886]    = ( l_42 [2918]);
assign l_41[2887]    = ( l_42 [2919]);
assign l_41[2888]    = ( l_42 [2920]);
assign l_41[2889]    = ( l_42 [2921]);
assign l_41[2890]    = ( l_42 [2922]);
assign l_41[2891]    = ( l_42 [2923]);
assign l_41[2892]    = ( l_42 [2924]);
assign l_41[2893]    = ( l_42 [2925]);
assign l_41[2894]    = ( l_42 [2926]);
assign l_41[2895]    = ( l_42 [2927]);
assign l_41[2896]    = ( l_42 [2928]);
assign l_41[2897]    = ( l_42 [2929]);
assign l_41[2898]    = ( l_42 [2930]);
assign l_41[2899]    = ( l_42 [2931]);
assign l_41[2900]    = ( l_42 [2932]);
assign l_41[2901]    = ( l_42 [2933]);
assign l_41[2902]    = ( l_42 [2934]);
assign l_41[2903]    = ( l_42 [2935]);
assign l_41[2904]    = ( l_42 [2936]);
assign l_41[2905]    = ( l_42 [2937]);
assign l_41[2906]    = ( l_42 [2938]);
assign l_41[2907]    = ( l_42 [2939]);
assign l_41[2908]    = ( l_42 [2940]);
assign l_41[2909]    = ( l_42 [2941]);
assign l_41[2910]    = ( l_42 [2942]);
assign l_41[2911]    = ( l_42 [2943]);
assign l_41[2912]    = ( l_42 [2944]);
assign l_41[2913]    = ( l_42 [2945]);
assign l_41[2914]    = ( l_42 [2946]);
assign l_41[2915]    = ( l_42 [2947]);
assign l_41[2916]    = ( l_42 [2948]);
assign l_41[2917]    = ( l_42 [2949]);
assign l_41[2918]    = ( l_42 [2950]);
assign l_41[2919]    = ( l_42 [2951]);
assign l_41[2920]    = ( l_42 [2952]);
assign l_41[2921]    = ( l_42 [2953]);
assign l_41[2922]    = ( l_42 [2954]);
assign l_41[2923]    = ( l_42 [2955]);
assign l_41[2924]    = ( l_42 [2956]);
assign l_41[2925]    = ( l_42 [2957]);
assign l_41[2926]    = ( l_42 [2958]);
assign l_41[2927]    = ( l_42 [2959]);
assign l_41[2928]    = ( l_42 [2960]);
assign l_41[2929]    = ( l_42 [2961]);
assign l_41[2930]    = ( l_42 [2962]);
assign l_41[2931]    = ( l_42 [2963]);
assign l_41[2932]    = ( l_42 [2964]);
assign l_41[2933]    = ( l_42 [2965]);
assign l_41[2934]    = ( l_42 [2966]);
assign l_41[2935]    = ( l_42 [2967]);
assign l_41[2936]    = ( l_42 [2968]);
assign l_41[2937]    = ( l_42 [2969]);
assign l_41[2938]    = ( l_42 [2970]);
assign l_41[2939]    = ( l_42 [2971]);
assign l_41[2940]    = ( l_42 [2972]);
assign l_41[2941]    = ( l_42 [2973]);
assign l_41[2942]    = ( l_42 [2974]);
assign l_41[2943]    = ( l_42 [2975]);
assign l_41[2944]    = ( l_42 [2976]);
assign l_41[2945]    = ( l_42 [2977]);
assign l_41[2946]    = ( l_42 [2978]);
assign l_41[2947]    = ( l_42 [2979]);
assign l_41[2948]    = ( l_42 [2980]);
assign l_41[2949]    = ( l_42 [2981]);
assign l_41[2950]    = ( l_42 [2982]);
assign l_41[2951]    = ( l_42 [2983]);
assign l_41[2952]    = ( l_42 [2984]);
assign l_41[2953]    = ( l_42 [2985]);
assign l_41[2954]    = ( l_42 [2986]);
assign l_41[2955]    = ( l_42 [2987]);
assign l_41[2956]    = ( l_42 [2988]);
assign l_41[2957]    = ( l_42 [2989]);
assign l_41[2958]    = ( l_42 [2990]);
assign l_41[2959]    = ( l_42 [2991]);
assign l_41[2960]    = ( l_42 [2992]);
assign l_41[2961]    = ( l_42 [2993]);
assign l_41[2962]    = ( l_42 [2994]);
assign l_41[2963]    = ( l_42 [2995]);
assign l_41[2964]    = ( l_42 [2996]);
assign l_41[2965]    = ( l_42 [2997]);
assign l_41[2966]    = ( l_42 [2998]);
assign l_41[2967]    = ( l_42 [2999]);
assign l_41[2968]    = ( l_42 [3000]);
assign l_41[2969]    = ( l_42 [3001]);
assign l_41[2970]    = ( l_42 [3002]);
assign l_41[2971]    = ( l_42 [3003]);
assign l_41[2972]    = ( l_42 [3004]);
assign l_41[2973]    = ( l_42 [3005]);
assign l_41[2974]    = ( l_42 [3006]);
assign l_41[2975]    = ( l_42 [3007]);
assign l_41[2976]    = ( l_42 [3008]);
assign l_41[2977]    = ( l_42 [3009]);
assign l_41[2978]    = ( l_42 [3010]);
assign l_41[2979]    = ( l_42 [3011]);
assign l_41[2980]    = ( l_42 [3012]);
assign l_41[2981]    = ( l_42 [3013]);
assign l_41[2982]    = ( l_42 [3014]);
assign l_41[2983]    = ( l_42 [3015]);
assign l_41[2984]    = ( l_42 [3016]);
assign l_41[2985]    = ( l_42 [3017]);
assign l_41[2986]    = ( l_42 [3018]);
assign l_41[2987]    = ( l_42 [3019]);
assign l_41[2988]    = ( l_42 [3020]);
assign l_41[2989]    = ( l_42 [3021]);
assign l_41[2990]    = ( l_42 [3022]);
assign l_41[2991]    = ( l_42 [3023]);
assign l_41[2992]    = ( l_42 [3024]);
assign l_41[2993]    = ( l_42 [3025]);
assign l_41[2994]    = ( l_42 [3026]);
assign l_41[2995]    = ( l_42 [3027]);
assign l_41[2996]    = ( l_42 [3028]);
assign l_41[2997]    = ( l_42 [3029]);
assign l_41[2998]    = ( l_42 [3030]);
assign l_41[2999]    = ( l_42 [3031]);
assign l_41[3000]    = ( l_42 [3032]);
assign l_41[3001]    = ( l_42 [3033]);
assign l_41[3002]    = ( l_42 [3034]);
assign l_41[3003]    = ( l_42 [3035]);
assign l_41[3004]    = ( l_42 [3036]);
assign l_41[3005]    = ( l_42 [3037]);
assign l_41[3006]    = ( l_42 [3038]);
assign l_41[3007]    = ( l_42 [3039]);
assign l_41[3008]    = ( l_42 [3040]);
assign l_41[3009]    = ( l_42 [3041]);
assign l_41[3010]    = ( l_42 [3042]);
assign l_41[3011]    = ( l_42 [3043]);
assign l_41[3012]    = ( l_42 [3044]);
assign l_41[3013]    = ( l_42 [3045]);
assign l_41[3014]    = ( l_42 [3046]);
assign l_41[3015]    = ( l_42 [3047]);
assign l_41[3016]    = ( l_42 [3048]);
assign l_41[3017]    = ( l_42 [3049]);
assign l_41[3018]    = ( l_42 [3050]);
assign l_41[3019]    = ( l_42 [3051]);
assign l_41[3020]    = ( l_42 [3052]);
assign l_41[3021]    = ( l_42 [3053]);
assign l_41[3022]    = ( l_42 [3054]);
assign l_41[3023]    = ( l_42 [3055]);
assign l_41[3024]    = ( l_42 [3056]);
assign l_41[3025]    = ( l_42 [3057]);
assign l_41[3026]    = ( l_42 [3058]);
assign l_41[3027]    = ( l_42 [3059]);
assign l_41[3028]    = ( l_42 [3060]);
assign l_41[3029]    = ( l_42 [3061]);
assign l_41[3030]    = ( l_42 [3062]);
assign l_41[3031]    = ( l_42 [3063]);
assign l_41[3032]    = ( l_42 [3064]);
assign l_41[3033]    = ( l_42 [3065]);
assign l_41[3034]    = ( l_42 [3066]);
assign l_41[3035]    = ( l_42 [3067]);
assign l_41[3036]    = ( l_42 [3068]);
assign l_41[3037]    = ( l_42 [3069]);
assign l_41[3038]    = ( l_42 [3070]);
assign l_41[3039]    = ( l_42 [3071]);
assign l_41[3040]    = ( l_42 [3072]);
assign l_41[3041]    = ( l_42 [3073]);
assign l_41[3042]    = ( l_42 [3074]);
assign l_41[3043]    = ( l_42 [3075]);
assign l_41[3044]    = ( l_42 [3076]);
assign l_41[3045]    = ( l_42 [3077]);
assign l_41[3046]    = ( l_42 [3078]);
assign l_41[3047]    = ( l_42 [3079]);
assign l_41[3048]    = ( l_42 [3080]);
assign l_41[3049]    = ( l_42 [3081]);
assign l_41[3050]    = ( l_42 [3082]);
assign l_41[3051]    = ( l_42 [3083]);
assign l_41[3052]    = ( l_42 [3084]);
assign l_41[3053]    = ( l_42 [3085]);
assign l_41[3054]    = ( l_42 [3086]);
assign l_41[3055]    = ( l_42 [3087]);
assign l_41[3056]    = ( l_42 [3088]);
assign l_41[3057]    = ( l_42 [3089]);
assign l_41[3058]    = ( l_42 [3090]);
assign l_41[3059]    = ( l_42 [3091]);
assign l_41[3060]    = ( l_42 [3092]);
assign l_41[3061]    = ( l_42 [3093]);
assign l_41[3062]    = ( l_42 [3094]);
assign l_41[3063]    = ( l_42 [3095]);
assign l_41[3064]    = ( l_42 [3096]);
assign l_41[3065]    = ( l_42 [3097]);
assign l_41[3066]    = ( l_42 [3098]);
assign l_41[3067]    = ( l_42 [3099]);
assign l_41[3068]    = ( l_42 [3100]);
assign l_41[3069]    = ( l_42 [3101]);
assign l_41[3070]    = ( l_42 [3102]);
assign l_41[3071]    = ( l_42 [3103]);
assign l_41[3072]    = ( l_42 [3104]);
assign l_41[3073]    = ( l_42 [3105]);
assign l_41[3074]    = ( l_42 [3106]);
assign l_41[3075]    = ( l_42 [3107]);
assign l_41[3076]    = ( l_42 [3108]);
assign l_41[3077]    = ( l_42 [3109]);
assign l_41[3078]    = ( l_42 [3110]);
assign l_41[3079]    = ( l_42 [3111]);
assign l_41[3080]    = ( l_42 [3112]);
assign l_41[3081]    = ( l_42 [3113]);
assign l_41[3082]    = ( l_42 [3114]);
assign l_41[3083]    = ( l_42 [3115]);
assign l_41[3084]    = ( l_42 [3116]);
assign l_41[3085]    = ( l_42 [3117]);
assign l_41[3086]    = ( l_42 [3118]);
assign l_41[3087]    = ( l_42 [3119]);
assign l_41[3088]    = ( l_42 [3120]);
assign l_41[3089]    = ( l_42 [3121]);
assign l_41[3090]    = ( l_42 [3122]);
assign l_41[3091]    = ( l_42 [3123]);
assign l_41[3092]    = ( l_42 [3124]);
assign l_41[3093]    = ( l_42 [3125]);
assign l_41[3094]    = ( l_42 [3126]);
assign l_41[3095]    = ( l_42 [3127]);
assign l_41[3096]    = ( l_42 [3128]);
assign l_41[3097]    = ( l_42 [3129]);
assign l_41[3098]    = ( l_42 [3130]);
assign l_41[3099]    = ( l_42 [3131]);
assign l_41[3100]    = ( l_42 [3132]);
assign l_41[3101]    = ( l_42 [3133]);
assign l_41[3102]    = ( l_42 [3134]);
assign l_41[3103]    = ( l_42 [3135]);
assign l_41[3104]    = ( l_42 [3136]);
assign l_41[3105]    = ( l_42 [3137]);
assign l_41[3106]    = ( l_42 [3138]);
assign l_41[3107]    = ( l_42 [3139]);
assign l_41[3108]    = ( l_42 [3140]);
assign l_41[3109]    = ( l_42 [3141]);
assign l_41[3110]    = ( l_42 [3142]);
assign l_41[3111]    = ( l_42 [3143]);
assign l_41[3112]    = ( l_42 [3144]);
assign l_41[3113]    = ( l_42 [3145]);
assign l_41[3114]    = ( l_42 [3146]);
assign l_41[3115]    = ( l_42 [3147]);
assign l_41[3116]    = ( l_42 [3148]);
assign l_41[3117]    = ( l_42 [3149]);
assign l_41[3118]    = ( l_42 [3150]);
assign l_41[3119]    = ( l_42 [3151]);
assign l_41[3120]    = ( l_42 [3152]);
assign l_41[3121]    = ( l_42 [3153]);
assign l_41[3122]    = ( l_42 [3154]);
assign l_41[3123]    = ( l_42 [3155]);
assign l_41[3124]    = ( l_42 [3156]);
assign l_41[3125]    = ( l_42 [3157]);
assign l_41[3126]    = ( l_42 [3158]);
assign l_41[3127]    = ( l_42 [3159]);
assign l_41[3128]    = ( l_42 [3160]);
assign l_41[3129]    = ( l_42 [3161]);
assign l_41[3130]    = ( l_42 [3162]);
assign l_41[3131]    = ( l_42 [3163]);
assign l_41[3132]    = ( l_42 [3164]);
assign l_41[3133]    = ( l_42 [3165]);
assign l_41[3134]    = ( l_42 [3166]);
assign l_41[3135]    = ( l_42 [3167]);
assign l_41[3136]    = ( l_42 [3168]);
assign l_41[3137]    = ( l_42 [3169]);
assign l_41[3138]    = ( l_42 [3170]);
assign l_41[3139]    = ( l_42 [3171]);
assign l_41[3140]    = ( l_42 [3172]);
assign l_41[3141]    = ( l_42 [3173]);
assign l_41[3142]    = ( l_42 [3174]);
assign l_41[3143]    = ( l_42 [3175]);
assign l_41[3144]    = ( l_42 [3176]);
assign l_41[3145]    = ( l_42 [3177]);
assign l_41[3146]    = ( l_42 [3178]);
assign l_41[3147]    = ( l_42 [3179]);
assign l_41[3148]    = ( l_42 [3180]);
assign l_41[3149]    = ( l_42 [3181]);
assign l_41[3150]    = ( l_42 [3182]);
assign l_41[3151]    = ( l_42 [3183]);
assign l_41[3152]    = ( l_42 [3184]);
assign l_41[3153]    = ( l_42 [3185]);
assign l_41[3154]    = ( l_42 [3186]);
assign l_41[3155]    = ( l_42 [3187]);
assign l_41[3156]    = ( l_42 [3188]);
assign l_41[3157]    = ( l_42 [3189]);
assign l_41[3158]    = ( l_42 [3190]);
assign l_41[3159]    = ( l_42 [3191]);
assign l_41[3160]    = ( l_42 [3192]);
assign l_41[3161]    = ( l_42 [3193]);
assign l_41[3162]    = ( l_42 [3194]);
assign l_41[3163]    = ( l_42 [3195]);
assign l_41[3164]    = ( l_42 [3196]);
assign l_41[3165]    = ( l_42 [3197]);
assign l_41[3166]    = ( l_42 [3198]);
assign l_41[3167]    = ( l_42 [3199]);
assign l_41[3168]    = ( l_42 [3200]);
assign l_41[3169]    = ( l_42 [3201]);
assign l_41[3170]    = ( l_42 [3202]);
assign l_41[3171]    = ( l_42 [3203]);
assign l_41[3172]    = ( l_42 [3204]);
assign l_41[3173]    = ( l_42 [3205]);
assign l_41[3174]    = ( l_42 [3206]);
assign l_41[3175]    = ( l_42 [3207]);
assign l_41[3176]    = ( l_42 [3208]);
assign l_41[3177]    = ( l_42 [3209]);
assign l_41[3178]    = ( l_42 [3210]);
assign l_41[3179]    = ( l_42 [3211]);
assign l_41[3180]    = ( l_42 [3212]);
assign l_41[3181]    = ( l_42 [3213]);
assign l_41[3182]    = ( l_42 [3214]);
assign l_41[3183]    = ( l_42 [3215]);
assign l_41[3184]    = ( l_42 [3216]);
assign l_41[3185]    = ( l_42 [3217]);
assign l_41[3186]    = ( l_42 [3218]);
assign l_41[3187]    = ( l_42 [3219]);
assign l_41[3188]    = ( l_42 [3220]);
assign l_41[3189]    = ( l_42 [3221]);
assign l_41[3190]    = ( l_42 [3222]);
assign l_41[3191]    = ( l_42 [3223]);
assign l_41[3192]    = ( l_42 [3224]);
assign l_41[3193]    = ( l_42 [3225]);
assign l_41[3194]    = ( l_42 [3226]);
assign l_41[3195]    = ( l_42 [3227]);
assign l_41[3196]    = ( l_42 [3228]);
assign l_41[3197]    = ( l_42 [3229]);
assign l_41[3198]    = ( l_42 [3230]);
assign l_41[3199]    = ( l_42 [3231]);
assign l_41[3200]    = ( l_42 [3232]);
assign l_41[3201]    = ( l_42 [3233]);
assign l_41[3202]    = ( l_42 [3234]);
assign l_41[3203]    = ( l_42 [3235]);
assign l_41[3204]    = ( l_42 [3236]);
assign l_41[3205]    = ( l_42 [3237]);
assign l_41[3206]    = ( l_42 [3238]);
assign l_41[3207]    = ( l_42 [3239]);
assign l_41[3208]    = ( l_42 [3240]);
assign l_41[3209]    = ( l_42 [3241]);
assign l_41[3210]    = ( l_42 [3242]);
assign l_41[3211]    = ( l_42 [3243]);
assign l_41[3212]    = ( l_42 [3244]);
assign l_41[3213]    = ( l_42 [3245]);
assign l_41[3214]    = ( l_42 [3246]);
assign l_41[3215]    = ( l_42 [3247]);
assign l_41[3216]    = ( l_42 [3248]);
assign l_41[3217]    = ( l_42 [3249]);
assign l_41[3218]    = ( l_42 [3250]);
assign l_41[3219]    = ( l_42 [3251]);
assign l_41[3220]    = ( l_42 [3252]);
assign l_41[3221]    = ( l_42 [3253]);
assign l_41[3222]    = ( l_42 [3254]);
assign l_41[3223]    = ( l_42 [3255]);
assign l_41[3224]    = ( l_42 [3256]);
assign l_41[3225]    = ( l_42 [3257]);
assign l_41[3226]    = ( l_42 [3258]);
assign l_41[3227]    = ( l_42 [3259]);
assign l_41[3228]    = ( l_42 [3260]);
assign l_41[3229]    = ( l_42 [3261]);
assign l_41[3230]    = ( l_42 [3262]);
assign l_41[3231]    = ( l_42 [3263]);
assign l_41[3232]    = ( l_42 [3264]);
assign l_41[3233]    = ( l_42 [3265]);
assign l_41[3234]    = ( l_42 [3266]);
assign l_41[3235]    = ( l_42 [3267]);
assign l_41[3236]    = ( l_42 [3268]);
assign l_41[3237]    = ( l_42 [3269]);
assign l_41[3238]    = ( l_42 [3270]);
assign l_41[3239]    = ( l_42 [3271]);
assign l_41[3240]    = ( l_42 [3272]);
assign l_41[3241]    = ( l_42 [3273]);
assign l_41[3242]    = ( l_42 [3274]);
assign l_41[3243]    = ( l_42 [3275]);
assign l_41[3244]    = ( l_42 [3276]);
assign l_41[3245]    = ( l_42 [3277]);
assign l_41[3246]    = ( l_42 [3278]);
assign l_41[3247]    = ( l_42 [3279]);
assign l_41[3248]    = ( l_42 [3280]);
assign l_41[3249]    = ( l_42 [3281]);
assign l_41[3250]    = ( l_42 [3282]);
assign l_41[3251]    = ( l_42 [3283]);
assign l_41[3252]    = ( l_42 [3284]);
assign l_41[3253]    = ( l_42 [3285]);
assign l_41[3254]    = ( l_42 [3286]);
assign l_41[3255]    = ( l_42 [3287]);
assign l_41[3256]    = ( l_42 [3288]);
assign l_41[3257]    = ( l_42 [3289]);
assign l_41[3258]    = ( l_42 [3290]);
assign l_41[3259]    = ( l_42 [3291]);
assign l_41[3260]    = ( l_42 [3292]);
assign l_41[3261]    = ( l_42 [3293]);
assign l_41[3262]    = ( l_42 [3294]);
assign l_41[3263]    = ( l_42 [3295]);
assign l_41[3264]    = ( l_42 [3296]);
assign l_41[3265]    = ( l_42 [3297]);
assign l_41[3266]    = ( l_42 [3298]);
assign l_41[3267]    = ( l_42 [3299]);
assign l_41[3268]    = ( l_42 [3300]);
assign l_41[3269]    = ( l_42 [3301]);
assign l_41[3270]    = ( l_42 [3302]);
assign l_41[3271]    = ( l_42 [3303]);
assign l_41[3272]    = ( l_42 [3304]);
assign l_41[3273]    = ( l_42 [3305]);
assign l_41[3274]    = ( l_42 [3306]);
assign l_41[3275]    = ( l_42 [3307]);
assign l_41[3276]    = ( l_42 [3308]);
assign l_41[3277]    = ( l_42 [3309]);
assign l_41[3278]    = ( l_42 [3310]);
assign l_41[3279]    = ( l_42 [3311]);
assign l_41[3280]    = ( l_42 [3312]);
assign l_41[3281]    = ( l_42 [3313]);
assign l_41[3282]    = ( l_42 [3314]);
assign l_41[3283]    = ( l_42 [3315]);
assign l_41[3284]    = ( l_42 [3316]);
assign l_41[3285]    = ( l_42 [3317]);
assign l_41[3286]    = ( l_42 [3318]);
assign l_41[3287]    = ( l_42 [3319]);
assign l_41[3288]    = ( l_42 [3320]);
assign l_41[3289]    = ( l_42 [3321]);
assign l_41[3290]    = ( l_42 [3322]);
assign l_41[3291]    = ( l_42 [3323]);
assign l_41[3292]    = ( l_42 [3324]);
assign l_41[3293]    = ( l_42 [3325]);
assign l_41[3294]    = ( l_42 [3326]);
assign l_41[3295]    = ( l_42 [3327]);
assign l_41[3296]    = ( l_42 [3328]);
assign l_41[3297]    = ( l_42 [3329]);
assign l_41[3298]    = ( l_42 [3330]);
assign l_41[3299]    = ( l_42 [3331]);
assign l_41[3300]    = ( l_42 [3332]);
assign l_41[3301]    = ( l_42 [3333]);
assign l_41[3302]    = ( l_42 [3334]);
assign l_41[3303]    = ( l_42 [3335]);
assign l_41[3304]    = ( l_42 [3336]);
assign l_41[3305]    = ( l_42 [3337]);
assign l_41[3306]    = ( l_42 [3338]);
assign l_41[3307]    = ( l_42 [3339]);
assign l_41[3308]    = ( l_42 [3340]);
assign l_41[3309]    = ( l_42 [3341]);
assign l_41[3310]    = ( l_42 [3342]);
assign l_41[3311]    = ( l_42 [3343]);
assign l_41[3312]    = ( l_42 [3344]);
assign l_41[3313]    = ( l_42 [3345]);
assign l_41[3314]    = ( l_42 [3346]);
assign l_41[3315]    = ( l_42 [3347]);
assign l_41[3316]    = ( l_42 [3348]);
assign l_41[3317]    = ( l_42 [3349]);
assign l_41[3318]    = ( l_42 [3350]);
assign l_41[3319]    = ( l_42 [3351]);
assign l_41[3320]    = ( l_42 [3352]);
assign l_41[3321]    = ( l_42 [3353]);
assign l_41[3322]    = ( l_42 [3354]);
assign l_41[3323]    = ( l_42 [3355]);
assign l_41[3324]    = ( l_42 [3356]);
assign l_41[3325]    = ( l_42 [3357]);
assign l_41[3326]    = ( l_42 [3358]);
assign l_41[3327]    = ( l_42 [3359]);
assign l_41[3328]    = ( l_42 [3360]);
assign l_41[3329]    = ( l_42 [3361]);
assign l_41[3330]    = ( l_42 [3362]);
assign l_41[3331]    = ( l_42 [3363]);
assign l_41[3332]    = ( l_42 [3364]);
assign l_41[3333]    = ( l_42 [3365]);
assign l_41[3334]    = ( l_42 [3366]);
assign l_41[3335]    = ( l_42 [3367]);
assign l_41[3336]    = ( l_42 [3368]);
assign l_41[3337]    = ( l_42 [3369]);
assign l_41[3338]    = ( l_42 [3370]);
assign l_41[3339]    = ( l_42 [3371]);
assign l_41[3340]    = ( l_42 [3372]);
assign l_41[3341]    = ( l_42 [3373]);
assign l_41[3342]    = ( l_42 [3374]);
assign l_41[3343]    = ( l_42 [3375]);
assign l_41[3344]    = ( l_42 [3376]);
assign l_41[3345]    = ( l_42 [3377]);
assign l_41[3346]    = ( l_42 [3378]);
assign l_41[3347]    = ( l_42 [3379]);
assign l_41[3348]    = ( l_42 [3380]);
assign l_41[3349]    = ( l_42 [3381]);
assign l_41[3350]    = ( l_42 [3382]);
assign l_41[3351]    = ( l_42 [3383]);
assign l_41[3352]    = ( l_42 [3384]);
assign l_41[3353]    = ( l_42 [3385]);
assign l_41[3354]    = ( l_42 [3386]);
assign l_41[3355]    = ( l_42 [3387]);
assign l_41[3356]    = ( l_42 [3388]);
assign l_41[3357]    = ( l_42 [3389]);
assign l_41[3358]    = ( l_42 [3390]);
assign l_41[3359]    = ( l_42 [3391]);
assign l_41[3360]    = ( l_42 [3392]);
assign l_41[3361]    = ( l_42 [3393]);
assign l_41[3362]    = ( l_42 [3394]);
assign l_41[3363]    = ( l_42 [3395]);
assign l_41[3364]    = ( l_42 [3396]);
assign l_41[3365]    = ( l_42 [3397]);
assign l_41[3366]    = ( l_42 [3398]);
assign l_41[3367]    = ( l_42 [3399]);
assign l_41[3368]    = ( l_42 [3400]);
assign l_41[3369]    = ( l_42 [3401]);
assign l_41[3370]    = ( l_42 [3402]);
assign l_41[3371]    = ( l_42 [3403]);
assign l_41[3372]    = ( l_42 [3404]);
assign l_41[3373]    = ( l_42 [3405]);
assign l_41[3374]    = ( l_42 [3406]);
assign l_41[3375]    = ( l_42 [3407]);
assign l_41[3376]    = ( l_42 [3408]);
assign l_41[3377]    = ( l_42 [3409]);
assign l_41[3378]    = ( l_42 [3410]);
assign l_41[3379]    = ( l_42 [3411]);
assign l_41[3380]    = ( l_42 [3412]);
assign l_41[3381]    = ( l_42 [3413]);
assign l_41[3382]    = ( l_42 [3414]);
assign l_41[3383]    = ( l_42 [3415]);
assign l_41[3384]    = ( l_42 [3416]);
assign l_41[3385]    = ( l_42 [3417]);
assign l_41[3386]    = ( l_42 [3418]);
assign l_41[3387]    = ( l_42 [3419]);
assign l_41[3388]    = ( l_42 [3420]);
assign l_41[3389]    = ( l_42 [3421]);
assign l_41[3390]    = ( l_42 [3422]);
assign l_41[3391]    = ( l_42 [3423]);
assign l_41[3392]    = ( l_42 [3424]);
assign l_41[3393]    = ( l_42 [3425]);
assign l_41[3394]    = ( l_42 [3426]);
assign l_41[3395]    = ( l_42 [3427]);
assign l_41[3396]    = ( l_42 [3428]);
assign l_41[3397]    = ( l_42 [3429]);
assign l_41[3398]    = ( l_42 [3430]);
assign l_41[3399]    = ( l_42 [3431]);
assign l_41[3400]    = ( l_42 [3432]);
assign l_41[3401]    = ( l_42 [3433]);
assign l_41[3402]    = ( l_42 [3434]);
assign l_41[3403]    = ( l_42 [3435]);
assign l_41[3404]    = ( l_42 [3436]);
assign l_41[3405]    = ( l_42 [3437]);
assign l_41[3406]    = ( l_42 [3438]);
assign l_41[3407]    = ( l_42 [3439]);
assign l_41[3408]    = ( l_42 [3440]);
assign l_41[3409]    = ( l_42 [3441]);
assign l_41[3410]    = ( l_42 [3442]);
assign l_41[3411]    = ( l_42 [3443]);
assign l_41[3412]    = ( l_42 [3444]);
assign l_41[3413]    = ( l_42 [3445]);
assign l_41[3414]    = ( l_42 [3446]);
assign l_41[3415]    = ( l_42 [3447]);
assign l_41[3416]    = ( l_42 [3448]);
assign l_41[3417]    = ( l_42 [3449]);
assign l_41[3418]    = ( l_42 [3450]);
assign l_41[3419]    = ( l_42 [3451]);
assign l_41[3420]    = ( l_42 [3452]);
assign l_41[3421]    = ( l_42 [3453]);
assign l_41[3422]    = ( l_42 [3454]);
assign l_41[3423]    = ( l_42 [3455]);
assign l_41[3424]    = ( l_42 [3456]);
assign l_41[3425]    = ( l_42 [3457]);
assign l_41[3426]    = ( l_42 [3458]);
assign l_41[3427]    = ( l_42 [3459]);
assign l_41[3428]    = ( l_42 [3460]);
assign l_41[3429]    = ( l_42 [3461]);
assign l_41[3430]    = ( l_42 [3462]);
assign l_41[3431]    = ( l_42 [3463]);
assign l_41[3432]    = ( l_42 [3464]);
assign l_41[3433]    = ( l_42 [3465]);
assign l_41[3434]    = ( l_42 [3466]);
assign l_41[3435]    = ( l_42 [3467]);
assign l_41[3436]    = ( l_42 [3468]);
assign l_41[3437]    = ( l_42 [3469]);
assign l_41[3438]    = ( l_42 [3470]);
assign l_41[3439]    = ( l_42 [3471]);
assign l_41[3440]    = ( l_42 [3472]);
assign l_41[3441]    = ( l_42 [3473]);
assign l_41[3442]    = ( l_42 [3474]);
assign l_41[3443]    = ( l_42 [3475]);
assign l_41[3444]    = ( l_42 [3476]);
assign l_41[3445]    = ( l_42 [3477]);
assign l_41[3446]    = ( l_42 [3478]);
assign l_41[3447]    = ( l_42 [3479]);
assign l_41[3448]    = ( l_42 [3480]);
assign l_41[3449]    = ( l_42 [3481]);
assign l_41[3450]    = ( l_42 [3482]);
assign l_41[3451]    = ( l_42 [3483]);
assign l_41[3452]    = ( l_42 [3484]);
assign l_41[3453]    = ( l_42 [3485]);
assign l_41[3454]    = ( l_42 [3486]);
assign l_41[3455]    = ( l_42 [3487]);
assign l_41[3456]    = ( l_42 [3488]);
assign l_41[3457]    = ( l_42 [3489]);
assign l_41[3458]    = ( l_42 [3490]);
assign l_41[3459]    = ( l_42 [3491]);
assign l_41[3460]    = ( l_42 [3492]);
assign l_41[3461]    = ( l_42 [3493]);
assign l_41[3462]    = ( l_42 [3494]);
assign l_41[3463]    = ( l_42 [3495]);
assign l_41[3464]    = ( l_42 [3496]);
assign l_41[3465]    = ( l_42 [3497]);
assign l_41[3466]    = ( l_42 [3498]);
assign l_41[3467]    = ( l_42 [3499]);
assign l_41[3468]    = ( l_42 [3500]);
assign l_41[3469]    = ( l_42 [3501]);
assign l_41[3470]    = ( l_42 [3502]);
assign l_41[3471]    = ( l_42 [3503]);
assign l_41[3472]    = ( l_42 [3504]);
assign l_41[3473]    = ( l_42 [3505]);
assign l_41[3474]    = ( l_42 [3506]);
assign l_41[3475]    = ( l_42 [3507]);
assign l_41[3476]    = ( l_42 [3508]);
assign l_41[3477]    = ( l_42 [3509]);
assign l_41[3478]    = ( l_42 [3510]);
assign l_41[3479]    = ( l_42 [3511]);
assign l_41[3480]    = ( l_42 [3512]);
assign l_41[3481]    = ( l_42 [3513]);
assign l_41[3482]    = ( l_42 [3514]);
assign l_41[3483]    = ( l_42 [3515]);
assign l_41[3484]    = ( l_42 [3516]);
assign l_41[3485]    = ( l_42 [3517]);
assign l_41[3486]    = ( l_42 [3518]);
assign l_41[3487]    = ( l_42 [3519]);
assign l_41[3488]    = ( l_42 [3520]);
assign l_41[3489]    = ( l_42 [3521]);
assign l_41[3490]    = ( l_42 [3522]);
assign l_41[3491]    = ( l_42 [3523]);
assign l_41[3492]    = ( l_42 [3524]);
assign l_41[3493]    = ( l_42 [3525]);
assign l_41[3494]    = ( l_42 [3526]);
assign l_41[3495]    = ( l_42 [3527]);
assign l_41[3496]    = ( l_42 [3528]);
assign l_41[3497]    = ( l_42 [3529]);
assign l_41[3498]    = ( l_42 [3530]);
assign l_41[3499]    = ( l_42 [3531]);
assign l_41[3500]    = ( l_42 [3532]);
assign l_41[3501]    = ( l_42 [3533]);
assign l_41[3502]    = ( l_42 [3534]);
assign l_41[3503]    = ( l_42 [3535]);
assign l_41[3504]    = ( l_42 [3536]);
assign l_41[3505]    = ( l_42 [3537]);
assign l_41[3506]    = ( l_42 [3538]);
assign l_41[3507]    = ( l_42 [3539]);
assign l_41[3508]    = ( l_42 [3540]);
assign l_41[3509]    = ( l_42 [3541]);
assign l_41[3510]    = ( l_42 [3542]);
assign l_41[3511]    = ( l_42 [3543]);
assign l_41[3512]    = ( l_42 [3544]);
assign l_41[3513]    = ( l_42 [3545]);
assign l_41[3514]    = ( l_42 [3546]);
assign l_41[3515]    = ( l_42 [3547]);
assign l_41[3516]    = ( l_42 [3548]);
assign l_41[3517]    = ( l_42 [3549]);
assign l_41[3518]    = ( l_42 [3550]);
assign l_41[3519]    = ( l_42 [3551]);
assign l_41[3520]    = ( l_42 [3552]);
assign l_41[3521]    = ( l_42 [3553]);
assign l_41[3522]    = ( l_42 [3554]);
assign l_41[3523]    = ( l_42 [3555]);
assign l_41[3524]    = ( l_42 [3556]);
assign l_41[3525]    = ( l_42 [3557]);
assign l_41[3526]    = ( l_42 [3558]);
assign l_41[3527]    = ( l_42 [3559]);
assign l_41[3528]    = ( l_42 [3560]);
assign l_41[3529]    = ( l_42 [3561]);
assign l_41[3530]    = ( l_42 [3562]);
assign l_41[3531]    = ( l_42 [3563]);
assign l_41[3532]    = ( l_42 [3564]);
assign l_41[3533]    = ( l_42 [3565]);
assign l_41[3534]    = ( l_42 [3566]);
assign l_41[3535]    = ( l_42 [3567]);
assign l_41[3536]    = ( l_42 [3568]);
assign l_41[3537]    = ( l_42 [3569]);
assign l_41[3538]    = ( l_42 [3570]);
assign l_41[3539]    = ( l_42 [3571]);
assign l_41[3540]    = ( l_42 [3572]);
assign l_41[3541]    = ( l_42 [3573]);
assign l_41[3542]    = ( l_42 [3574]);
assign l_41[3543]    = ( l_42 [3575]);
assign l_41[3544]    = ( l_42 [3576]);
assign l_41[3545]    = ( l_42 [3577]);
assign l_41[3546]    = ( l_42 [3578]);
assign l_41[3547]    = ( l_42 [3579]);
assign l_41[3548]    = ( l_42 [3580]);
assign l_41[3549]    = ( l_42 [3581]);
assign l_41[3550]    = ( l_42 [3582]);
assign l_41[3551]    = ( l_42 [3583]);
assign l_41[3552]    = ( l_42 [3584]);
assign l_41[3553]    = ( l_42 [3585]);
assign l_41[3554]    = ( l_42 [3586]);
assign l_41[3555]    = ( l_42 [3587]);
assign l_41[3556]    = ( l_42 [3588]);
assign l_41[3557]    = ( l_42 [3589]);
assign l_41[3558]    = ( l_42 [3590]);
assign l_41[3559]    = ( l_42 [3591]);
assign l_41[3560]    = ( l_42 [3592]);
assign l_41[3561]    = ( l_42 [3593]);
assign l_41[3562]    = ( l_42 [3594]);
assign l_41[3563]    = ( l_42 [3595]);
assign l_41[3564]    = ( l_42 [3596]);
assign l_41[3565]    = ( l_42 [3597]);
assign l_41[3566]    = ( l_42 [3598]);
assign l_41[3567]    = ( l_42 [3599]);
assign l_41[3568]    = ( l_42 [3600]);
assign l_41[3569]    = ( l_42 [3601]);
assign l_41[3570]    = ( l_42 [3602]);
assign l_41[3571]    = ( l_42 [3603]);
assign l_41[3572]    = ( l_42 [3604]);
assign l_41[3573]    = ( l_42 [3605]);
assign l_41[3574]    = ( l_42 [3606]);
assign l_41[3575]    = ( l_42 [3607]);
assign l_41[3576]    = ( l_42 [3608]);
assign l_41[3577]    = ( l_42 [3609]);
assign l_41[3578]    = ( l_42 [3610]);
assign l_41[3579]    = ( l_42 [3611]);
assign l_41[3580]    = ( l_42 [3612]);
assign l_41[3581]    = ( l_42 [3613]);
assign l_41[3582]    = ( l_42 [3614]);
assign l_41[3583]    = ( l_42 [3615]);
assign l_41[3584]    = ( l_42 [3616]);
assign l_41[3585]    = ( l_42 [3617]);
assign l_41[3586]    = ( l_42 [3618]);
assign l_41[3587]    = ( l_42 [3619]);
assign l_41[3588]    = ( l_42 [3620]);
assign l_41[3589]    = ( l_42 [3621]);
assign l_41[3590]    = ( l_42 [3622]);
assign l_41[3591]    = ( l_42 [3623]);
assign l_41[3592]    = ( l_42 [3624]);
assign l_41[3593]    = ( l_42 [3625]);
assign l_41[3594]    = ( l_42 [3626]);
assign l_41[3595]    = ( l_42 [3627]);
assign l_41[3596]    = ( l_42 [3628]);
assign l_41[3597]    = ( l_42 [3629]);
assign l_41[3598]    = ( l_42 [3630]);
assign l_41[3599]    = ( l_42 [3631]);
assign l_41[3600]    = ( l_42 [3632]);
assign l_41[3601]    = ( l_42 [3633]);
assign l_41[3602]    = ( l_42 [3634]);
assign l_41[3603]    = ( l_42 [3635]);
assign l_41[3604]    = ( l_42 [3636]);
assign l_41[3605]    = ( l_42 [3637]);
assign l_41[3606]    = ( l_42 [3638]);
assign l_41[3607]    = ( l_42 [3639]);
assign l_41[3608]    = ( l_42 [3640]);
assign l_41[3609]    = ( l_42 [3641]);
assign l_41[3610]    = ( l_42 [3642]);
assign l_41[3611]    = ( l_42 [3643]);
assign l_41[3612]    = ( l_42 [3644]);
assign l_41[3613]    = ( l_42 [3645]);
assign l_41[3614]    = ( l_42 [3646]);
assign l_41[3615]    = ( l_42 [3647]);
assign l_41[3616]    = ( l_42 [3648]);
assign l_41[3617]    = ( l_42 [3649]);
assign l_41[3618]    = ( l_42 [3650]);
assign l_41[3619]    = ( l_42 [3651]);
assign l_41[3620]    = ( l_42 [3652]);
assign l_41[3621]    = ( l_42 [3653]);
assign l_41[3622]    = ( l_42 [3654]);
assign l_41[3623]    = ( l_42 [3655]);
assign l_41[3624]    = ( l_42 [3656]);
assign l_41[3625]    = ( l_42 [3657]);
assign l_41[3626]    = ( l_42 [3658]);
assign l_41[3627]    = ( l_42 [3659]);
assign l_41[3628]    = ( l_42 [3660]);
assign l_41[3629]    = ( l_42 [3661]);
assign l_41[3630]    = ( l_42 [3662]);
assign l_41[3631]    = ( l_42 [3663]);
assign l_41[3632]    = ( l_42 [3664]);
assign l_41[3633]    = ( l_42 [3665]);
assign l_41[3634]    = ( l_42 [3666]);
assign l_41[3635]    = ( l_42 [3667]);
assign l_41[3636]    = ( l_42 [3668]);
assign l_41[3637]    = ( l_42 [3669]);
assign l_41[3638]    = ( l_42 [3670]);
assign l_41[3639]    = ( l_42 [3671]);
assign l_41[3640]    = ( l_42 [3672]);
assign l_41[3641]    = ( l_42 [3673]);
assign l_41[3642]    = ( l_42 [3674]);
assign l_41[3643]    = ( l_42 [3675]);
assign l_41[3644]    = ( l_42 [3676]);
assign l_41[3645]    = ( l_42 [3677]);
assign l_41[3646]    = ( l_42 [3678]);
assign l_41[3647]    = ( l_42 [3679]);
assign l_41[3648]    = ( l_42 [3680]);
assign l_41[3649]    = ( l_42 [3681]);
assign l_41[3650]    = ( l_42 [3682]);
assign l_41[3651]    = ( l_42 [3683]);
assign l_41[3652]    = ( l_42 [3684]);
assign l_41[3653]    = ( l_42 [3685]);
assign l_41[3654]    = ( l_42 [3686]);
assign l_41[3655]    = ( l_42 [3687]);
assign l_41[3656]    = ( l_42 [3688]);
assign l_41[3657]    = ( l_42 [3689]);
assign l_41[3658]    = ( l_42 [3690]);
assign l_41[3659]    = ( l_42 [3691]);
assign l_41[3660]    = ( l_42 [3692]);
assign l_41[3661]    = ( l_42 [3693]);
assign l_41[3662]    = ( l_42 [3694]);
assign l_41[3663]    = ( l_42 [3695]);
assign l_41[3664]    = ( l_42 [3696]);
assign l_41[3665]    = ( l_42 [3697]);
assign l_41[3666]    = ( l_42 [3698]);
assign l_41[3667]    = ( l_42 [3699]);
assign l_41[3668]    = ( l_42 [3700]);
assign l_41[3669]    = ( l_42 [3701]);
assign l_41[3670]    = ( l_42 [3702]);
assign l_41[3671]    = ( l_42 [3703]);
assign l_41[3672]    = ( l_42 [3704]);
assign l_41[3673]    = ( l_42 [3705]);
assign l_41[3674]    = ( l_42 [3706]);
assign l_41[3675]    = ( l_42 [3707]);
assign l_41[3676]    = ( l_42 [3708]);
assign l_41[3677]    = ( l_42 [3709]);
assign l_41[3678]    = ( l_42 [3710]);
assign l_41[3679]    = ( l_42 [3711]);
assign l_41[3680]    = ( l_42 [3712]);
assign l_41[3681]    = ( l_42 [3713]);
assign l_41[3682]    = ( l_42 [3714]);
assign l_41[3683]    = ( l_42 [3715]);
assign l_41[3684]    = ( l_42 [3716]);
assign l_41[3685]    = ( l_42 [3717]);
assign l_41[3686]    = ( l_42 [3718]);
assign l_41[3687]    = ( l_42 [3719]);
assign l_41[3688]    = ( l_42 [3720]);
assign l_41[3689]    = ( l_42 [3721]);
assign l_41[3690]    = ( l_42 [3722]);
assign l_41[3691]    = ( l_42 [3723]);
assign l_41[3692]    = ( l_42 [3724]);
assign l_41[3693]    = ( l_42 [3725]);
assign l_41[3694]    = ( l_42 [3726]);
assign l_41[3695]    = ( l_42 [3727]);
assign l_41[3696]    = ( l_42 [3728]);
assign l_41[3697]    = ( l_42 [3729]);
assign l_41[3698]    = ( l_42 [3730]);
assign l_41[3699]    = ( l_42 [3731]);
assign l_41[3700]    = ( l_42 [3732]);
assign l_41[3701]    = ( l_42 [3733]);
assign l_41[3702]    = ( l_42 [3734]);
assign l_41[3703]    = ( l_42 [3735]);
assign l_41[3704]    = ( l_42 [3736]);
assign l_41[3705]    = ( l_42 [3737]);
assign l_41[3706]    = ( l_42 [3738]);
assign l_41[3707]    = ( l_42 [3739]);
assign l_41[3708]    = ( l_42 [3740]);
assign l_41[3709]    = ( l_42 [3741]);
assign l_41[3710]    = ( l_42 [3742]);
assign l_41[3711]    = ( l_42 [3743]);
assign l_41[3712]    = ( l_42 [3744]);
assign l_41[3713]    = ( l_42 [3745]);
assign l_41[3714]    = ( l_42 [3746]);
assign l_41[3715]    = ( l_42 [3747]);
assign l_41[3716]    = ( l_42 [3748]);
assign l_41[3717]    = ( l_42 [3749]);
assign l_41[3718]    = ( l_42 [3750]);
assign l_41[3719]    = ( l_42 [3751]);
assign l_41[3720]    = ( l_42 [3752]);
assign l_41[3721]    = ( l_42 [3753]);
assign l_41[3722]    = ( l_42 [3754]);
assign l_41[3723]    = ( l_42 [3755]);
assign l_41[3724]    = ( l_42 [3756]);
assign l_41[3725]    = ( l_42 [3757]);
assign l_41[3726]    = ( l_42 [3758]);
assign l_41[3727]    = ( l_42 [3759]);
assign l_41[3728]    = ( l_42 [3760]);
assign l_41[3729]    = ( l_42 [3761]);
assign l_41[3730]    = ( l_42 [3762]);
assign l_41[3731]    = ( l_42 [3763]);
assign l_41[3732]    = ( l_42 [3764]);
assign l_41[3733]    = ( l_42 [3765]);
assign l_41[3734]    = ( l_42 [3766]);
assign l_41[3735]    = ( l_42 [3767]);
assign l_41[3736]    = ( l_42 [3768]);
assign l_41[3737]    = ( l_42 [3769]);
assign l_41[3738]    = ( l_42 [3770]);
assign l_41[3739]    = ( l_42 [3771]);
assign l_41[3740]    = ( l_42 [3772]);
assign l_41[3741]    = ( l_42 [3773]);
assign l_41[3742]    = ( l_42 [3774]);
assign l_41[3743]    = ( l_42 [3775]);
assign l_41[3744]    = ( l_42 [3776]);
assign l_41[3745]    = ( l_42 [3777]);
assign l_41[3746]    = ( l_42 [3778]);
assign l_41[3747]    = ( l_42 [3779]);
assign l_41[3748]    = ( l_42 [3780]);
assign l_41[3749]    = ( l_42 [3781]);
assign l_41[3750]    = ( l_42 [3782]);
assign l_41[3751]    = ( l_42 [3783]);
assign l_41[3752]    = ( l_42 [3784]);
assign l_41[3753]    = ( l_42 [3785]);
assign l_41[3754]    = ( l_42 [3786]);
assign l_41[3755]    = ( l_42 [3787]);
assign l_41[3756]    = ( l_42 [3788]);
assign l_41[3757]    = ( l_42 [3789]);
assign l_41[3758]    = ( l_42 [3790]);
assign l_41[3759]    = ( l_42 [3791]);
assign l_41[3760]    = ( l_42 [3792]);
assign l_41[3761]    = ( l_42 [3793]);
assign l_41[3762]    = ( l_42 [3794]);
assign l_41[3763]    = ( l_42 [3795]);
assign l_41[3764]    = ( l_42 [3796]);
assign l_41[3765]    = ( l_42 [3797]);
assign l_41[3766]    = ( l_42 [3798]);
assign l_41[3767]    = ( l_42 [3799]);
assign l_41[3768]    = ( l_42 [3800]);
assign l_41[3769]    = ( l_42 [3801]);
assign l_41[3770]    = ( l_42 [3802]);
assign l_41[3771]    = ( l_42 [3803]);
assign l_41[3772]    = ( l_42 [3804]);
assign l_41[3773]    = ( l_42 [3805]);
assign l_41[3774]    = ( l_42 [3806]);
assign l_41[3775]    = ( l_42 [3807]);
assign l_41[3776]    = ( l_42 [3808]);
assign l_41[3777]    = ( l_42 [3809]);
assign l_41[3778]    = ( l_42 [3810]);
assign l_41[3779]    = ( l_42 [3811]);
assign l_41[3780]    = ( l_42 [3812]);
assign l_41[3781]    = ( l_42 [3813]);
assign l_41[3782]    = ( l_42 [3814]);
assign l_41[3783]    = ( l_42 [3815]);
assign l_41[3784]    = ( l_42 [3816]);
assign l_41[3785]    = ( l_42 [3817]);
assign l_41[3786]    = ( l_42 [3818]);
assign l_41[3787]    = ( l_42 [3819]);
assign l_41[3788]    = ( l_42 [3820]);
assign l_41[3789]    = ( l_42 [3821]);
assign l_41[3790]    = ( l_42 [3822]);
assign l_41[3791]    = ( l_42 [3823]);
assign l_41[3792]    = ( l_42 [3824]);
assign l_41[3793]    = ( l_42 [3825]);
assign l_41[3794]    = ( l_42 [3826]);
assign l_41[3795]    = ( l_42 [3827]);
assign l_41[3796]    = ( l_42 [3828]);
assign l_41[3797]    = ( l_42 [3829]);
assign l_41[3798]    = ( l_42 [3830]);
assign l_41[3799]    = ( l_42 [3831]);
assign l_41[3800]    = ( l_42 [3832]);
assign l_41[3801]    = ( l_42 [3833]);
assign l_41[3802]    = ( l_42 [3834]);
assign l_41[3803]    = ( l_42 [3835]);
assign l_41[3804]    = ( l_42 [3836]);
assign l_41[3805]    = ( l_42 [3837]);
assign l_41[3806]    = ( l_42 [3838]);
assign l_41[3807]    = ( l_42 [3839]);
assign l_41[3808]    = ( l_42 [3840]);
assign l_41[3809]    = ( l_42 [3841]);
assign l_41[3810]    = ( l_42 [3842]);
assign l_41[3811]    = ( l_42 [3843]);
assign l_41[3812]    = ( l_42 [3844]);
assign l_41[3813]    = ( l_42 [3845]);
assign l_41[3814]    = ( l_42 [3846]);
assign l_41[3815]    = ( l_42 [3847]);
assign l_41[3816]    = ( l_42 [3848]);
assign l_41[3817]    = ( l_42 [3849]);
assign l_41[3818]    = ( l_42 [3850]);
assign l_41[3819]    = ( l_42 [3851]);
assign l_41[3820]    = ( l_42 [3852]);
assign l_41[3821]    = ( l_42 [3853]);
assign l_41[3822]    = ( l_42 [3854]);
assign l_41[3823]    = ( l_42 [3855]);
assign l_41[3824]    = ( l_42 [3856]);
assign l_41[3825]    = ( l_42 [3857]);
assign l_41[3826]    = ( l_42 [3858]);
assign l_41[3827]    = ( l_42 [3859]);
assign l_41[3828]    = ( l_42 [3860]);
assign l_41[3829]    = ( l_42 [3861]);
assign l_41[3830]    = ( l_42 [3862]);
assign l_41[3831]    = ( l_42 [3863]);
assign l_41[3832]    = ( l_42 [3864]);
assign l_41[3833]    = ( l_42 [3865]);
assign l_41[3834]    = ( l_42 [3866]);
assign l_41[3835]    = ( l_42 [3867]);
assign l_41[3836]    = ( l_42 [3868]);
assign l_41[3837]    = ( l_42 [3869]);
assign l_41[3838]    = ( l_42 [3870]);
assign l_41[3839]    = ( l_42 [3871]);
assign l_41[3840]    = ( l_42 [3872]);
assign l_41[3841]    = ( l_42 [3873]);
assign l_41[3842]    = ( l_42 [3874]);
assign l_41[3843]    = ( l_42 [3875]);
assign l_41[3844]    = ( l_42 [3876]);
assign l_41[3845]    = ( l_42 [3877]);
assign l_41[3846]    = ( l_42 [3878]);
assign l_41[3847]    = ( l_42 [3879]);
assign l_41[3848]    = ( l_42 [3880]);
assign l_41[3849]    = ( l_42 [3881]);
assign l_41[3850]    = ( l_42 [3882]);
assign l_41[3851]    = ( l_42 [3883]);
assign l_41[3852]    = ( l_42 [3884]);
assign l_41[3853]    = ( l_42 [3885]);
assign l_41[3854]    = ( l_42 [3886]);
assign l_41[3855]    = ( l_42 [3887]);
assign l_41[3856]    = ( l_42 [3888]);
assign l_41[3857]    = ( l_42 [3889]);
assign l_41[3858]    = ( l_42 [3890]);
assign l_41[3859]    = ( l_42 [3891]);
assign l_41[3860]    = ( l_42 [3892]);
assign l_41[3861]    = ( l_42 [3893]);
assign l_41[3862]    = ( l_42 [3894]);
assign l_41[3863]    = ( l_42 [3895]);
assign l_41[3864]    = ( l_42 [3896]);
assign l_41[3865]    = ( l_42 [3897]);
assign l_41[3866]    = ( l_42 [3898]);
assign l_41[3867]    = ( l_42 [3899]);
assign l_41[3868]    = ( l_42 [3900]);
assign l_41[3869]    = ( l_42 [3901]);
assign l_41[3870]    = ( l_42 [3902]);
assign l_41[3871]    = ( l_42 [3903]);
assign l_41[3872]    = ( l_42 [3904]);
assign l_41[3873]    = ( l_42 [3905]);
assign l_41[3874]    = ( l_42 [3906]);
assign l_41[3875]    = ( l_42 [3907]);
assign l_41[3876]    = ( l_42 [3908]);
assign l_41[3877]    = ( l_42 [3909]);
assign l_41[3878]    = ( l_42 [3910]);
assign l_41[3879]    = ( l_42 [3911]);
assign l_41[3880]    = ( l_42 [3912]);
assign l_41[3881]    = ( l_42 [3913]);
assign l_41[3882]    = ( l_42 [3914]);
assign l_41[3883]    = ( l_42 [3915]);
assign l_41[3884]    = ( l_42 [3916]);
assign l_41[3885]    = ( l_42 [3917]);
assign l_41[3886]    = ( l_42 [3918]);
assign l_41[3887]    = ( l_42 [3919]);
assign l_41[3888]    = ( l_42 [3920]);
assign l_41[3889]    = ( l_42 [3921]);
assign l_41[3890]    = ( l_42 [3922]);
assign l_41[3891]    = ( l_42 [3923]);
assign l_41[3892]    = ( l_42 [3924]);
assign l_41[3893]    = ( l_42 [3925]);
assign l_41[3894]    = ( l_42 [3926]);
assign l_41[3895]    = ( l_42 [3927]);
assign l_41[3896]    = ( l_42 [3928]);
assign l_41[3897]    = ( l_42 [3929]);
assign l_41[3898]    = ( l_42 [3930]);
assign l_41[3899]    = ( l_42 [3931]);
assign l_41[3900]    = ( l_42 [3932]);
assign l_41[3901]    = ( l_42 [3933]);
assign l_41[3902]    = ( l_42 [3934]);
assign l_41[3903]    = ( l_42 [3935]);
assign l_41[3904]    = ( l_42 [3936]);
assign l_41[3905]    = ( l_42 [3937]);
assign l_41[3906]    = ( l_42 [3938]);
assign l_41[3907]    = ( l_42 [3939]);
assign l_41[3908]    = ( l_42 [3940]);
assign l_41[3909]    = ( l_42 [3941]);
assign l_41[3910]    = ( l_42 [3942]);
assign l_41[3911]    = ( l_42 [3943]);
assign l_41[3912]    = ( l_42 [3944]);
assign l_41[3913]    = ( l_42 [3945]);
assign l_41[3914]    = ( l_42 [3946]);
assign l_41[3915]    = ( l_42 [3947]);
assign l_41[3916]    = ( l_42 [3948]);
assign l_41[3917]    = ( l_42 [3949]);
assign l_41[3918]    = ( l_42 [3950]);
assign l_41[3919]    = ( l_42 [3951]);
assign l_41[3920]    = ( l_42 [3952]);
assign l_41[3921]    = ( l_42 [3953]);
assign l_41[3922]    = ( l_42 [3954]);
assign l_41[3923]    = ( l_42 [3955]);
assign l_41[3924]    = ( l_42 [3956]);
assign l_41[3925]    = ( l_42 [3957]);
assign l_41[3926]    = ( l_42 [3958]);
assign l_41[3927]    = ( l_42 [3959]);
assign l_41[3928]    = ( l_42 [3960]);
assign l_41[3929]    = ( l_42 [3961]);
assign l_41[3930]    = ( l_42 [3962]);
assign l_41[3931]    = ( l_42 [3963]);
assign l_41[3932]    = ( l_42 [3964]);
assign l_41[3933]    = ( l_42 [3965]);
assign l_41[3934]    = ( l_42 [3966]);
assign l_41[3935]    = ( l_42 [3967]);
assign l_41[3936]    = ( l_42 [3968]);
assign l_41[3937]    = ( l_42 [3969]);
assign l_41[3938]    = ( l_42 [3970]);
assign l_41[3939]    = ( l_42 [3971]);
assign l_41[3940]    = ( l_42 [3972]);
assign l_41[3941]    = ( l_42 [3973]);
assign l_41[3942]    = ( l_42 [3974]);
assign l_41[3943]    = ( l_42 [3975]);
assign l_41[3944]    = ( l_42 [3976]);
assign l_41[3945]    = ( l_42 [3977]);
assign l_41[3946]    = ( l_42 [3978]);
assign l_41[3947]    = ( l_42 [3979]);
assign l_41[3948]    = ( l_42 [3980]);
assign l_41[3949]    = ( l_42 [3981]);
assign l_41[3950]    = ( l_42 [3982]);
assign l_41[3951]    = ( l_42 [3983]);
assign l_41[3952]    = ( l_42 [3984]);
assign l_41[3953]    = ( l_42 [3985]);
assign l_41[3954]    = ( l_42 [3986]);
assign l_41[3955]    = ( l_42 [3987]);
assign l_41[3956]    = ( l_42 [3988]);
assign l_41[3957]    = ( l_42 [3989]);
assign l_41[3958]    = ( l_42 [3990]);
assign l_41[3959]    = ( l_42 [3991]);
assign l_41[3960]    = ( l_42 [3992]);
assign l_41[3961]    = ( l_42 [3993]);
assign l_41[3962]    = ( l_42 [3994]);
assign l_41[3963]    = ( l_42 [3995]);
assign l_41[3964]    = ( l_42 [3996]);
assign l_41[3965]    = ( l_42 [3997]);
assign l_41[3966]    = ( l_42 [3998]);
assign l_41[3967]    = ( l_42 [3999]);
assign l_41[3968]    = ( l_42 [4000]);
assign l_41[3969]    = ( l_42 [4001]);
assign l_41[3970]    = ( l_42 [4002]);
assign l_41[3971]    = ( l_42 [4003]);
assign l_41[3972]    = ( l_42 [4004]);
assign l_41[3973]    = ( l_42 [4005]);
assign l_41[3974]    = ( l_42 [4006]);
assign l_41[3975]    = ( l_42 [4007]);
assign l_41[3976]    = ( l_42 [4008]);
assign l_41[3977]    = ( l_42 [4009]);
assign l_41[3978]    = ( l_42 [4010]);
assign l_41[3979]    = ( l_42 [4011]);
assign l_41[3980]    = ( l_42 [4012]);
assign l_41[3981]    = ( l_42 [4013]);
assign l_41[3982]    = ( l_42 [4014]);
assign l_41[3983]    = ( l_42 [4015]);
assign l_41[3984]    = ( l_42 [4016]);
assign l_41[3985]    = ( l_42 [4017]);
assign l_41[3986]    = ( l_42 [4018]);
assign l_41[3987]    = ( l_42 [4019]);
assign l_41[3988]    = ( l_42 [4020]);
assign l_41[3989]    = ( l_42 [4021]);
assign l_41[3990]    = ( l_42 [4022]);
assign l_41[3991]    = ( l_42 [4023]);
assign l_41[3992]    = ( l_42 [4024]);
assign l_41[3993]    = ( l_42 [4025]);
assign l_41[3994]    = ( l_42 [4026]);
assign l_41[3995]    = ( l_42 [4027]);
assign l_41[3996]    = ( l_42 [4028]);
assign l_41[3997]    = ( l_42 [4029]);
assign l_41[3998]    = ( l_42 [4030]);
assign l_41[3999]    = ( l_42 [4031]);
assign l_41[4000]    = ( l_42 [4032]);
assign l_41[4001]    = ( l_42 [4033]);
assign l_41[4002]    = ( l_42 [4034]);
assign l_41[4003]    = ( l_42 [4035]);
assign l_41[4004]    = ( l_42 [4036]);
assign l_41[4005]    = ( l_42 [4037]);
assign l_41[4006]    = ( l_42 [4038]);
assign l_41[4007]    = ( l_42 [4039]);
assign l_41[4008]    = ( l_42 [4040]);
assign l_41[4009]    = ( l_42 [4041]);
assign l_41[4010]    = ( l_42 [4042]);
assign l_41[4011]    = ( l_42 [4043]);
assign l_41[4012]    = ( l_42 [4044]);
assign l_41[4013]    = ( l_42 [4045]);
assign l_41[4014]    = ( l_42 [4046]);
assign l_41[4015]    = ( l_42 [4047]);
assign l_41[4016]    = ( l_42 [4048]);
assign l_41[4017]    = ( l_42 [4049]);
assign l_41[4018]    = ( l_42 [4050]);
assign l_41[4019]    = ( l_42 [4051]);
assign l_41[4020]    = ( l_42 [4052]);
assign l_41[4021]    = ( l_42 [4053]);
assign l_41[4022]    = ( l_42 [4054]);
assign l_41[4023]    = ( l_42 [4055]);
assign l_41[4024]    = ( l_42 [4056]);
assign l_41[4025]    = ( l_42 [4057]);
assign l_41[4026]    = ( l_42 [4058]);
assign l_41[4027]    = ( l_42 [4059]);
assign l_41[4028]    = ( l_42 [4060]);
assign l_41[4029]    = ( l_42 [4061]);
assign l_41[4030]    = ( l_42 [4062]);
assign l_41[4031]    = ( l_42 [4063]);
assign l_41[4032]    = ( l_42 [4064]);
assign l_41[4033]    = ( l_42 [4065]);
assign l_41[4034]    = ( l_42 [4066]);
assign l_41[4035]    = ( l_42 [4067]);
assign l_41[4036]    = ( l_42 [4068]);
assign l_41[4037]    = ( l_42 [4069]);
assign l_41[4038]    = ( l_42 [4070]);
assign l_41[4039]    = ( l_42 [4071]);
assign l_41[4040]    = ( l_42 [4072]);
assign l_41[4041]    = ( l_42 [4073]);
assign l_41[4042]    = ( l_42 [4074]);
assign l_41[4043]    = ( l_42 [4075]);
assign l_41[4044]    = ( l_42 [4076]);
assign l_41[4045]    = ( l_42 [4077]);
assign l_41[4046]    = ( l_42 [4078]);
assign l_41[4047]    = ( l_42 [4079]);
assign l_41[4048]    = ( l_42 [4080]);
assign l_41[4049]    = ( l_42 [4081]);
assign l_41[4050]    = ( l_42 [4082]);
assign l_41[4051]    = ( l_42 [4083]);
assign l_41[4052]    = ( l_42 [4084]);
assign l_41[4053]    = ( l_42 [4085]);
assign l_41[4054]    = ( l_42 [4086]);
assign l_41[4055]    = ( l_42 [4087]);
assign l_41[4056]    = ( l_42 [4088]);
assign l_41[4057]    = ( l_42 [4089]);
assign l_41[4058]    = ( l_42 [4090]);
assign l_41[4059]    = ( l_42 [4091]);
assign l_41[4060]    = ( l_42 [4092]);
assign l_41[4061]    = ( l_42 [4093]);
assign l_41[4062]    = ( l_42 [4094]);
assign l_41[4063]    = ( l_42 [4095]);
assign l_41[4064]    = ( l_42 [4096]);
assign l_41[4065]    = ( l_42 [4097]);
assign l_41[4066]    = ( l_42 [4098]);
assign l_41[4067]    = ( l_42 [4099]);
assign l_41[4068]    = ( l_42 [4100]);
assign l_41[4069]    = ( l_42 [4101]);
assign l_41[4070]    = ( l_42 [4102]);
assign l_41[4071]    = ( l_42 [4103]);
assign l_41[4072]    = ( l_42 [4104]);
assign l_41[4073]    = ( l_42 [4105]);
assign l_41[4074]    = ( l_42 [4106]);
assign l_41[4075]    = ( l_42 [4107]);
assign l_41[4076]    = ( l_42 [4108]);
assign l_41[4077]    = ( l_42 [4109]);
assign l_41[4078]    = ( l_42 [4110]);
assign l_41[4079]    = ( l_42 [4111]);
assign l_41[4080]    = ( l_42 [4112]);
assign l_41[4081]    = ( l_42 [4113]);
assign l_41[4082]    = ( l_42 [4114]);
assign l_41[4083]    = ( l_42 [4115]);
assign l_41[4084]    = ( l_42 [4116]);
assign l_41[4085]    = ( l_42 [4117]);
assign l_41[4086]    = ( l_42 [4118]);
assign l_41[4087]    = ( l_42 [4119]);
assign l_41[4088]    = ( l_42 [4120]);
assign l_41[4089]    = ( l_42 [4121]);
assign l_41[4090]    = ( l_42 [4122]);
assign l_41[4091]    = ( l_42 [4123]);
assign l_41[4092]    = ( l_42 [4124]);
assign l_41[4093]    = ( l_42 [4125]);
assign l_41[4094]    = ( l_42 [4126]);
assign l_41[4095]    = ( l_42 [4127]);
assign l_41[4096]    = ( l_42 [4128]);
assign l_41[4097]    = ( l_42 [4129]);
assign l_41[4098]    = ( l_42 [4130]);
assign l_41[4099]    = ( l_42 [4131]);
assign l_41[4100]    = ( l_42 [4132]);
assign l_41[4101]    = ( l_42 [4133]);
assign l_41[4102]    = ( l_42 [4134]);
assign l_41[4103]    = ( l_42 [4135]);
assign l_41[4104]    = ( l_42 [4136]);
assign l_41[4105]    = ( l_42 [4137]);
assign l_41[4106]    = ( l_42 [4138]);
assign l_41[4107]    = ( l_42 [4139]);
assign l_41[4108]    = ( l_42 [4140]);
assign l_41[4109]    = ( l_42 [4141]);
assign l_41[4110]    = ( l_42 [4142]);
assign l_41[4111]    = ( l_42 [4143]);
assign l_41[4112]    = ( l_42 [4144]);
assign l_41[4113]    = ( l_42 [4145]);
assign l_41[4114]    = ( l_42 [4146]);
assign l_41[4115]    = ( l_42 [4147]);
assign l_41[4116]    = ( l_42 [4148]);
assign l_41[4117]    = ( l_42 [4149]);
assign l_41[4118]    = ( l_42 [4150]);
assign l_41[4119]    = ( l_42 [4151]);
assign l_41[4120]    = ( l_42 [4152]);
assign l_41[4121]    = ( l_42 [4153]);
assign l_41[4122]    = ( l_42 [4154]);
assign l_41[4123]    = ( l_42 [4155]);
assign l_41[4124]    = ( l_42 [4156]);
assign l_41[4125]    = ( l_42 [4157]);
assign l_41[4126]    = ( l_42 [4158]);
assign l_41[4127]    = ( l_42 [4159]);
assign l_41[4128]    = ( l_42 [4160]);
assign l_41[4129]    = ( l_42 [4161]);
assign l_41[4130]    = ( l_42 [4162] & !i[1820]) | ( l_42 [4163] &  i[1820]);
assign l_41[4131]    = ( l_42 [4164] & !i[1820]) | ( l_42 [4165] &  i[1820]);
assign l_41[4132]    = ( l_42 [4166] & !i[1820]) | ( l_42 [4167] &  i[1820]);
assign l_41[4133]    = ( l_42 [4168] & !i[1820]) | ( l_42 [4169] &  i[1820]);
assign l_41[4134]    = ( l_42 [4170] & !i[1820]) | ( l_42 [4171] &  i[1820]);
assign l_41[4135]    = ( l_42 [4172] & !i[1820]) | ( l_42 [4173] &  i[1820]);
assign l_41[4136]    = ( l_42 [4174] & !i[1820]) | ( l_42 [4175] &  i[1820]);
assign l_41[4137]    = ( l_42 [4176] & !i[1820]) | ( l_42 [4177] &  i[1820]);
assign l_41[4138]    = ( l_42 [4178] & !i[1820]) | ( l_42 [4179] &  i[1820]);
assign l_41[4139]    = ( l_42 [4180] & !i[1820]) | ( l_42 [4181] &  i[1820]);
assign l_41[4140]    = ( l_42 [4182] & !i[1820]) | ( l_42 [4183] &  i[1820]);
assign l_41[4141]    = ( l_42 [4184] & !i[1820]) | ( l_42 [4185] &  i[1820]);
assign l_41[4142]    = ( l_42 [4186] & !i[1820]) | ( l_42 [4187] &  i[1820]);
assign l_41[4143]    = ( l_42 [4188] & !i[1820]) | ( l_42 [4189] &  i[1820]);
assign l_41[4144]    = ( l_42 [4190] & !i[1820]) | ( l_42 [4191] &  i[1820]);
assign l_41[4145]    = ( l_42 [4192] & !i[1820]) | ( l_42 [4193] &  i[1820]);
assign l_41[4146]    = ( l_42 [4194] & !i[1820]) | ( l_42 [4195] &  i[1820]);
assign l_41[4147]    = ( l_42 [4196] & !i[1820]) | ( l_42 [4197] &  i[1820]);
assign l_41[4148]    = ( l_42 [4198] & !i[1820]) | ( l_42 [4199] &  i[1820]);
assign l_41[4149]    = ( l_42 [4200] & !i[1820]) | ( l_42 [4201] &  i[1820]);
assign l_41[4150]    = ( l_42 [4202] & !i[1820]) | ( l_42 [4203] &  i[1820]);
assign l_41[4151]    = ( l_42 [4204] & !i[1820]) | ( l_42 [4205] &  i[1820]);
assign l_41[4152]    = ( l_42 [4206] & !i[1820]) | ( l_42 [4207] &  i[1820]);
assign l_41[4153]    = ( l_42 [4208] & !i[1820]) | ( l_42 [4209] &  i[1820]);
assign l_41[4154]    = ( l_42 [4210] & !i[1820]) | ( l_42 [4211] &  i[1820]);
assign l_41[4155]    = ( l_42 [4212] & !i[1820]) | ( l_42 [4213] &  i[1820]);
assign l_41[4156]    = ( l_42 [4214] & !i[1820]) | ( l_42 [4215] &  i[1820]);
assign l_41[4157]    = ( l_42 [4216] & !i[1820]) | ( l_42 [4217] &  i[1820]);
assign l_41[4158]    = ( l_42 [4218] & !i[1820]) | ( l_42 [4219] &  i[1820]);
assign l_41[4159]    = ( l_42 [4220] & !i[1820]) | ( l_42 [4221] &  i[1820]);
assign l_41[4160]    = ( l_42 [4222] & !i[1820]) | ( l_42 [4223] &  i[1820]);
assign l_41[4161]    = ( l_42 [4224] & !i[1820]) | ( l_42 [4225] &  i[1820]);
assign l_41[4162]    = ( l_42 [4226] & !i[1820]) | ( l_42 [4227] &  i[1820]);
assign l_41[4163]    = ( l_42 [4228] & !i[1820]) | ( l_42 [4229] &  i[1820]);
assign l_41[4164]    = ( l_42 [4230] & !i[1820]) | ( l_42 [4231] &  i[1820]);
assign l_41[4165]    = ( l_42 [4232] & !i[1820]) | ( l_42 [4233] &  i[1820]);
assign l_41[4166]    = ( l_42 [4234] & !i[1820]) | ( l_42 [4235] &  i[1820]);
assign l_41[4167]    = ( l_42 [4236] & !i[1820]) | ( l_42 [4237] &  i[1820]);
assign l_41[4168]    = ( l_42 [4238] & !i[1820]) | ( l_42 [4239] &  i[1820]);
assign l_41[4169]    = ( l_42 [4240] & !i[1820]) | ( l_42 [4241] &  i[1820]);
assign l_41[4170]    = ( l_42 [4242] & !i[1820]) | ( l_42 [4243] &  i[1820]);
assign l_41[4171]    = ( l_42 [4244] & !i[1820]) | ( l_42 [4245] &  i[1820]);
assign l_41[4172]    = ( l_42 [4246] & !i[1820]) | ( l_42 [4247] &  i[1820]);
assign l_41[4173]    = ( l_42 [4248] & !i[1820]) | ( l_42 [4249] &  i[1820]);
assign l_41[4174]    = ( l_42 [4250] & !i[1820]) | ( l_42 [4251] &  i[1820]);
assign l_41[4175]    = ( l_42 [4252] & !i[1820]) | ( l_42 [4253] &  i[1820]);
assign l_41[4176]    = ( l_42 [4254] & !i[1820]) | ( l_42 [4255] &  i[1820]);
assign l_41[4177]    = ( l_42 [4256] & !i[1820]) | ( l_42 [4257] &  i[1820]);
assign l_41[4178]    = ( l_42 [4258] & !i[1820]) | ( l_42 [4259] &  i[1820]);
assign l_41[4179]    = ( l_42 [4260] & !i[1820]) | ( l_42 [4261] &  i[1820]);
assign l_41[4180]    = ( l_42 [4262] & !i[1820]) | ( l_42 [4263] &  i[1820]);
assign l_41[4181]    = ( l_42 [4264] & !i[1820]) | ( l_42 [4265] &  i[1820]);
assign l_41[4182]    = ( l_42 [4266] & !i[1820]) | ( l_42 [4267] &  i[1820]);
assign l_41[4183]    = ( l_42 [4268] & !i[1820]) | ( l_42 [4269] &  i[1820]);
assign l_41[4184]    = ( l_42 [4270] & !i[1820]) | ( l_42 [4271] &  i[1820]);
assign l_41[4185]    = ( l_42 [4272] & !i[1820]) | ( l_42 [4273] &  i[1820]);
assign l_41[4186]    = ( l_42 [4274] & !i[1820]) | ( l_42 [4275] &  i[1820]);
assign l_41[4187]    = ( l_42 [4276] & !i[1820]) | ( l_42 [4277] &  i[1820]);
assign l_41[4188]    = ( l_42 [4278] & !i[1820]) | ( l_42 [4279] &  i[1820]);
assign l_41[4189]    = ( l_42 [4280] & !i[1820]) | ( l_42 [4281] &  i[1820]);
assign l_41[4190]    = ( l_42 [4282] & !i[1820]) | ( l_42 [4283] &  i[1820]);
assign l_41[4191]    = ( l_42 [4284] & !i[1820]) | ( l_42 [4285] &  i[1820]);
assign l_41[4192]    = ( l_42 [4286] & !i[1820]) | ( l_42 [4287] &  i[1820]);
assign l_41[4193]    = ( l_42 [4288] & !i[1820]) | ( l_42 [4289] &  i[1820]);
assign l_41[4194]    = ( l_42 [4290] & !i[1820]) | ( l_42 [4291] &  i[1820]);
assign l_41[4195]    = ( l_42 [4292] & !i[1820]) | ( l_42 [4293] &  i[1820]);
assign l_41[4196]    = ( l_42 [4294] & !i[1820]) | ( l_42 [4295] &  i[1820]);
assign l_41[4197]    = ( l_42 [4296] & !i[1820]) | ( l_42 [4297] &  i[1820]);
assign l_41[4198]    = ( l_42 [4298] & !i[1820]) | ( l_42 [4299] &  i[1820]);
assign l_41[4199]    = ( l_42 [4300] & !i[1820]) | ( l_42 [4301] &  i[1820]);
assign l_41[4200]    = ( l_42 [4302] & !i[1820]) | ( l_42 [4303] &  i[1820]);
assign l_41[4201]    = ( l_42 [4304] & !i[1820]) | ( l_42 [4305] &  i[1820]);
assign l_41[4202]    = ( l_42 [4306] & !i[1820]) | ( l_42 [4307] &  i[1820]);
assign l_41[4203]    = ( l_42 [4308] & !i[1820]) | ( l_42 [4309] &  i[1820]);
assign l_41[4204]    = ( l_42 [4310] & !i[1820]) | ( l_42 [4311] &  i[1820]);
assign l_41[4205]    = ( l_42 [4312] & !i[1820]) | ( l_42 [4313] &  i[1820]);
assign l_41[4206]    = ( l_42 [4314] & !i[1820]) | ( l_42 [4315] &  i[1820]);
assign l_41[4207]    = ( l_42 [4316] & !i[1820]) | ( l_42 [4317] &  i[1820]);
assign l_41[4208]    = ( l_42 [4318] & !i[1820]) | ( l_42 [4319] &  i[1820]);
assign l_41[4209]    = ( l_42 [4320] & !i[1820]) | ( l_42 [4321] &  i[1820]);
assign l_41[4210]    = ( l_42 [4322] & !i[1820]) | ( l_42 [4323] &  i[1820]);
assign l_41[4211]    = ( l_42 [4324] & !i[1820]) | ( l_42 [4325] &  i[1820]);
assign l_41[4212]    = ( l_42 [4326] & !i[1820]) | ( l_42 [4327] &  i[1820]);
assign l_41[4213]    = ( l_42 [4328] & !i[1820]) | ( l_42 [4329] &  i[1820]);
assign l_41[4214]    = ( l_42 [4330] & !i[1820]) | ( l_42 [4331] &  i[1820]);
assign l_41[4215]    = ( l_42 [4332] & !i[1820]) | ( l_42 [4333] &  i[1820]);
assign l_41[4216]    = ( l_42 [4334] & !i[1820]) | ( l_42 [4335] &  i[1820]);
assign l_41[4217]    = ( l_42 [4336] & !i[1820]) | ( l_42 [4337] &  i[1820]);
assign l_41[4218]    = ( l_42 [4338] & !i[1820]) | ( l_42 [4339] &  i[1820]);
assign l_41[4219]    = ( l_42 [4340] & !i[1820]) | ( l_42 [4341] &  i[1820]);
assign l_41[4220]    = ( l_42 [4342] & !i[1820]) | ( l_42 [4343] &  i[1820]);
assign l_41[4221]    = ( l_42 [4344] & !i[1820]) | ( l_42 [4345] &  i[1820]);
assign l_41[4222]    = ( l_42 [4346] & !i[1820]) | ( l_42 [4347] &  i[1820]);
assign l_41[4223]    = ( l_42 [4348] & !i[1820]) | ( l_42 [4349] &  i[1820]);
assign l_41[4224]    = ( l_42 [4350] & !i[1820]) | ( l_42 [4351] &  i[1820]);
assign l_41[4225]    = ( l_42 [4352] & !i[1820]) | ( l_42 [4353] &  i[1820]);
assign l_41[4226]    = ( l_42 [4354] & !i[1820]) | ( l_42 [4355] &  i[1820]);
assign l_41[4227]    = ( l_42 [4356] & !i[1820]) | ( l_42 [4357] &  i[1820]);
assign l_41[4228]    = ( l_42 [4358] & !i[1820]) | ( l_42 [4359] &  i[1820]);
assign l_41[4229]    = ( l_42 [4360] & !i[1820]) | ( l_42 [4361] &  i[1820]);
assign l_41[4230]    = ( l_42 [4362] & !i[1820]) | ( l_42 [4363] &  i[1820]);
assign l_41[4231]    = ( l_42 [4364] & !i[1820]) | ( l_42 [4365] &  i[1820]);
assign l_41[4232]    = ( l_42 [4366] & !i[1820]) | ( l_42 [4367] &  i[1820]);
assign l_41[4233]    = ( l_42 [4368] & !i[1820]) | ( l_42 [4369] &  i[1820]);
assign l_41[4234]    = ( l_42 [4370] & !i[1820]) | ( l_42 [4371] &  i[1820]);
assign l_41[4235]    = ( l_42 [4372] & !i[1820]) | ( l_42 [4373] &  i[1820]);
assign l_41[4236]    = ( l_42 [4374] & !i[1820]) | ( l_42 [4375] &  i[1820]);
assign l_41[4237]    = ( l_42 [4376] & !i[1820]) | ( l_42 [4377] &  i[1820]);
assign l_41[4238]    = ( l_42 [4378] & !i[1820]) | ( l_42 [4379] &  i[1820]);
assign l_41[4239]    = ( l_42 [4380] & !i[1820]) | ( l_42 [4381] &  i[1820]);
assign l_41[4240]    = ( l_42 [4382] & !i[1820]) | ( l_42 [4383] &  i[1820]);
assign l_41[4241]    = ( l_42 [4384] & !i[1820]) | ( l_42 [4385] &  i[1820]);
assign l_41[4242]    = ( l_42 [4386] & !i[1820]) | ( l_42 [4387] &  i[1820]);
assign l_41[4243]    = ( l_42 [4388] & !i[1820]) | ( l_42 [4389] &  i[1820]);
assign l_41[4244]    = ( l_42 [4390] & !i[1820]) | ( l_42 [4391] &  i[1820]);
assign l_41[4245]    = ( l_42 [4392] & !i[1820]) | ( l_42 [4393] &  i[1820]);
assign l_41[4246]    = ( l_42 [4394] & !i[1820]) | ( l_42 [4395] &  i[1820]);
assign l_41[4247]    = ( l_42 [4396] & !i[1820]) | ( l_42 [4397] &  i[1820]);
assign l_41[4248]    = ( l_42 [4398] & !i[1820]) | ( l_42 [4399] &  i[1820]);
assign l_41[4249]    = ( l_42 [4400] & !i[1820]) | ( l_42 [4401] &  i[1820]);
assign l_41[4250]    = ( l_42 [4402] & !i[1820]) | ( l_42 [4403] &  i[1820]);
assign l_41[4251]    = ( l_42 [4404] & !i[1820]) | ( l_42 [4405] &  i[1820]);
assign l_41[4252]    = ( l_42 [4406] & !i[1820]) | ( l_42 [4407] &  i[1820]);
assign l_41[4253]    = ( l_42 [4408] & !i[1820]) | ( l_42 [4409] &  i[1820]);
assign l_41[4254]    = ( l_42 [4410] & !i[1820]) | ( l_42 [4411] &  i[1820]);
assign l_41[4255]    = ( l_42 [4412] & !i[1820]) | ( l_42 [4413] &  i[1820]);
assign l_41[4256]    = ( l_42 [4414] & !i[1820]) | ( l_42 [4415] &  i[1820]);
assign l_41[4257]    = ( l_42 [4416] & !i[1820]) | ( l_42 [4417] &  i[1820]);
assign l_41[4258]    = ( l_42 [4418] & !i[1820]) | ( l_42 [4419] &  i[1820]);
assign l_41[4259]    = ( l_42 [4420] & !i[1820]) | ( l_42 [4421] &  i[1820]);
assign l_41[4260]    = ( l_42 [4422] & !i[1820]) | ( l_42 [4423] &  i[1820]);
assign l_41[4261]    = ( l_42 [4424] & !i[1820]) | ( l_42 [4425] &  i[1820]);
assign l_41[4262]    = ( l_42 [4426] & !i[1820]) | ( l_42 [4427] &  i[1820]);
assign l_41[4263]    = ( l_42 [4428] & !i[1820]) | ( l_42 [4429] &  i[1820]);
assign l_41[4264]    = ( l_42 [4430] & !i[1820]) | ( l_42 [4431] &  i[1820]);
assign l_41[4265]    = ( l_42 [4432] & !i[1820]) | ( l_42 [4433] &  i[1820]);
assign l_41[4266]    = ( l_42 [4434] & !i[1820]) | ( l_42 [4435] &  i[1820]);
assign l_41[4267]    = ( l_42 [4436] & !i[1820]) | ( l_42 [4437] &  i[1820]);
assign l_41[4268]    = ( l_42 [4438] & !i[1820]) | ( l_42 [4439] &  i[1820]);
assign l_41[4269]    = ( l_42 [4440] & !i[1820]) | ( l_42 [4441] &  i[1820]);
assign l_41[4270]    = ( l_42 [4442] & !i[1820]) | ( l_42 [4443] &  i[1820]);
assign l_41[4271]    = ( l_42 [4444] & !i[1820]) | ( l_42 [4445] &  i[1820]);
assign l_41[4272]    = ( l_42 [4446] & !i[1820]) | ( l_42 [4447] &  i[1820]);
assign l_41[4273]    = ( l_42 [4448] & !i[1820]) | ( l_42 [4449] &  i[1820]);
assign l_41[4274]    = ( l_42 [4450] & !i[1820]) | ( l_42 [4451] &  i[1820]);
assign l_41[4275]    = ( l_42 [4452] & !i[1820]) | ( l_42 [4453] &  i[1820]);
assign l_41[4276]    = ( l_42 [4454] & !i[1820]) | ( l_42 [4455] &  i[1820]);
assign l_41[4277]    = ( l_42 [4456] & !i[1820]) | ( l_42 [4457] &  i[1820]);
assign l_41[4278]    = ( l_42 [4458] & !i[1820]) | ( l_42 [4459] &  i[1820]);
assign l_41[4279]    = ( l_42 [4460] & !i[1820]) | ( l_42 [4461] &  i[1820]);
assign l_41[4280]    = ( l_42 [4462] & !i[1820]) | ( l_42 [4463] &  i[1820]);
assign l_41[4281]    = ( l_42 [4464] & !i[1820]) | ( l_42 [4465] &  i[1820]);
assign l_41[4282]    = ( l_42 [4466] & !i[1820]) | ( l_42 [4467] &  i[1820]);
assign l_41[4283]    = ( l_42 [4468] & !i[1820]) | ( l_42 [4469] &  i[1820]);
assign l_41[4284]    = ( l_42 [4470] & !i[1820]) | ( l_42 [4471] &  i[1820]);
assign l_41[4285]    = ( l_42 [4472] & !i[1820]) | ( l_42 [4473] &  i[1820]);
assign l_41[4286]    = ( l_42 [4474] & !i[1820]) | ( l_42 [4475] &  i[1820]);
assign l_41[4287]    = ( l_42 [4476] & !i[1820]) | ( l_42 [4477] &  i[1820]);
assign l_41[4288]    = ( l_42 [4478] & !i[1820]) | ( l_42 [4479] &  i[1820]);
assign l_41[4289]    = ( l_42 [4480] & !i[1820]) | ( l_42 [4481] &  i[1820]);
assign l_41[4290]    = ( l_42 [4482] & !i[1820]) | ( l_42 [4483] &  i[1820]);
assign l_41[4291]    = ( l_42 [4484] & !i[1820]) | ( l_42 [4485] &  i[1820]);
assign l_41[4292]    = ( l_42 [4486] & !i[1820]) | ( l_42 [4487] &  i[1820]);
assign l_41[4293]    = ( l_42 [4488] & !i[1820]) | ( l_42 [4489] &  i[1820]);
assign l_41[4294]    = ( l_42 [4490] & !i[1820]) | ( l_42 [4491] &  i[1820]);
assign l_41[4295]    = ( l_42 [4492] & !i[1820]) | ( l_42 [4493] &  i[1820]);
assign l_41[4296]    = ( l_42 [4494] & !i[1820]) | ( l_42 [4495] &  i[1820]);
assign l_41[4297]    = ( l_42 [4496] & !i[1820]) | ( l_42 [4497] &  i[1820]);
assign l_41[4298]    = ( l_42 [4498] & !i[1820]) | ( l_42 [4499] &  i[1820]);
assign l_41[4299]    = ( l_42 [4500] & !i[1820]) | ( l_42 [4501] &  i[1820]);
assign l_41[4300]    = ( l_42 [4502] & !i[1820]) | ( l_42 [4503] &  i[1820]);
assign l_41[4301]    = ( l_42 [4504] & !i[1820]) | ( l_42 [4505] &  i[1820]);
assign l_41[4302]    = ( l_42 [4506] & !i[1820]) | ( l_42 [4507] &  i[1820]);
assign l_41[4303]    = ( l_42 [4508] & !i[1820]) | ( l_42 [4509] &  i[1820]);
assign l_41[4304]    = ( l_42 [4510] & !i[1820]) | ( l_42 [4511] &  i[1820]);
assign l_41[4305]    = ( l_42 [4512] & !i[1820]) | ( l_42 [4513] &  i[1820]);
assign l_41[4306]    = ( l_42 [4514] & !i[1820]) | ( l_42 [4515] &  i[1820]);
assign l_41[4307]    = ( l_42 [4516] & !i[1820]) | ( l_42 [4517] &  i[1820]);
assign l_41[4308]    = ( l_42 [4518] & !i[1820]) | ( l_42 [4519] &  i[1820]);
assign l_41[4309]    = ( l_42 [4520] & !i[1820]) | ( l_42 [4521] &  i[1820]);
assign l_41[4310]    = ( l_42 [4522] & !i[1820]) | ( l_42 [4523] &  i[1820]);
assign l_41[4311]    = ( l_42 [4524] & !i[1820]) | ( l_42 [4525] &  i[1820]);
assign l_41[4312]    = ( l_42 [4526] & !i[1820]) | ( l_42 [4527] &  i[1820]);
assign l_41[4313]    = ( l_42 [4528] & !i[1820]) | ( l_42 [4529] &  i[1820]);
assign l_41[4314]    = ( l_42 [4530] & !i[1820]) | ( l_42 [4531] &  i[1820]);
assign l_41[4315]    = ( l_42 [4532] & !i[1820]) | ( l_42 [4533] &  i[1820]);
assign l_41[4316]    = ( l_42 [4534] & !i[1820]) | ( l_42 [4535] &  i[1820]);
assign l_41[4317]    = ( l_42 [4536] & !i[1820]) | ( l_42 [4537] &  i[1820]);
assign l_41[4318]    = ( l_42 [4538] & !i[1820]) | ( l_42 [4539] &  i[1820]);
assign l_41[4319]    = ( l_42 [4540] & !i[1820]) | ( l_42 [4541] &  i[1820]);
assign l_41[4320]    = ( l_42 [4542] & !i[1820]) | ( l_42 [4543] &  i[1820]);
assign l_41[4321]    = ( l_42 [4544] & !i[1820]) | ( l_42 [4545] &  i[1820]);
assign l_41[4322]    = ( l_42 [4546] & !i[1820]) | ( l_42 [4547] &  i[1820]);
assign l_41[4323]    = ( l_42 [4548] & !i[1820]) | ( l_42 [4549] &  i[1820]);
assign l_41[4324]    = ( l_42 [4550] & !i[1820]) | ( l_42 [4551] &  i[1820]);
assign l_41[4325]    = ( l_42 [4552] & !i[1820]) | ( l_42 [4553] &  i[1820]);
assign l_41[4326]    = ( l_42 [4554] & !i[1820]) | ( l_42 [4555] &  i[1820]);
assign l_41[4327]    = ( l_42 [4556] & !i[1820]) | ( l_42 [4557] &  i[1820]);
assign l_41[4328]    = ( l_42 [4558] & !i[1820]) | ( l_42 [4559] &  i[1820]);
assign l_41[4329]    = ( l_42 [4560] & !i[1820]) | ( l_42 [4561] &  i[1820]);
assign l_41[4330]    = ( l_42 [4562] & !i[1820]) | ( l_42 [4563] &  i[1820]);
assign l_41[4331]    = ( l_42 [4564] & !i[1820]) | ( l_42 [4565] &  i[1820]);
assign l_41[4332]    = ( l_42 [4566] & !i[1820]) | ( l_42 [4567] &  i[1820]);
assign l_41[4333]    = ( l_42 [4568] & !i[1820]) | ( l_42 [4569] &  i[1820]);
assign l_41[4334]    = ( l_42 [4570] & !i[1820]) | ( l_42 [4571] &  i[1820]);
assign l_41[4335]    = ( l_42 [4572] & !i[1820]) | ( l_42 [4573] &  i[1820]);
assign l_41[4336]    = ( l_42 [4574] & !i[1820]) | ( l_42 [4575] &  i[1820]);
assign l_41[4337]    = ( l_42 [4576] & !i[1820]) | ( l_42 [4577] &  i[1820]);
assign l_41[4338]    = ( l_42 [4578] & !i[1820]) | ( l_42 [4579] &  i[1820]);
assign l_41[4339]    = ( l_42 [4580] & !i[1820]) | ( l_42 [4581] &  i[1820]);
assign l_41[4340]    = ( l_42 [4582] & !i[1820]) | ( l_42 [4583] &  i[1820]);
assign l_41[4341]    = ( l_42 [4584] & !i[1820]) | ( l_42 [4585] &  i[1820]);
assign l_41[4342]    = ( l_42 [4586] & !i[1820]) | ( l_42 [4587] &  i[1820]);
assign l_41[4343]    = ( l_42 [4588] & !i[1820]) | ( l_42 [4589] &  i[1820]);
assign l_41[4344]    = ( l_42 [4590] & !i[1820]) | ( l_42 [4591] &  i[1820]);
assign l_41[4345]    = ( l_42 [4592] & !i[1820]) | ( l_42 [4593] &  i[1820]);
assign l_41[4346]    = ( l_42 [4594] & !i[1820]) | ( l_42 [4595] &  i[1820]);
assign l_41[4347]    = ( l_42 [4596] & !i[1820]) | ( l_42 [4597] &  i[1820]);
assign l_41[4348]    = ( l_42 [4598] & !i[1820]) | ( l_42 [4599] &  i[1820]);
assign l_41[4349]    = ( l_42 [4600] & !i[1820]) | ( l_42 [4601] &  i[1820]);
assign l_41[4350]    = ( l_42 [4602] & !i[1820]) | ( l_42 [4603] &  i[1820]);
assign l_41[4351]    = ( l_42 [4604] & !i[1820]) | ( l_42 [4605] &  i[1820]);
assign l_41[4352]    = ( l_42 [4606] & !i[1820]) | ( l_42 [4607] &  i[1820]);
assign l_41[4353]    = ( l_42 [4608] & !i[1820]) | ( l_42 [4609] &  i[1820]);
assign l_41[4354]    = ( l_42 [4610] & !i[1820]) | ( l_42 [4611] &  i[1820]);
assign l_41[4355]    = ( l_42 [4612] & !i[1820]) | ( l_42 [4613] &  i[1820]);
assign l_41[4356]    = ( l_42 [4614] & !i[1820]) | ( l_42 [4615] &  i[1820]);
assign l_41[4357]    = ( l_42 [4616] & !i[1820]) | ( l_42 [4617] &  i[1820]);
assign l_41[4358]    = ( l_42 [4618] & !i[1820]) | ( l_42 [4619] &  i[1820]);
assign l_41[4359]    = ( l_42 [4620] & !i[1820]) | ( l_42 [4621] &  i[1820]);
assign l_41[4360]    = ( l_42 [4622] & !i[1820]) | ( l_42 [4623] &  i[1820]);
assign l_41[4361]    = ( l_42 [4624] & !i[1820]) | ( l_42 [4625] &  i[1820]);
assign l_41[4362]    = ( l_42 [4626] & !i[1820]) | ( l_42 [4627] &  i[1820]);
assign l_41[4363]    = ( l_42 [4628] & !i[1820]) | ( l_42 [4629] &  i[1820]);
assign l_41[4364]    = ( l_42 [4630] & !i[1820]) | ( l_42 [4631] &  i[1820]);
assign l_41[4365]    = ( l_42 [4632] & !i[1820]) | ( l_42 [4633] &  i[1820]);
assign l_41[4366]    = ( l_42 [4634] & !i[1820]) | ( l_42 [4635] &  i[1820]);
assign l_41[4367]    = ( l_42 [4636] & !i[1820]) | ( l_42 [4637] &  i[1820]);
assign l_41[4368]    = ( l_42 [4638] & !i[1820]) | ( l_42 [4639] &  i[1820]);
assign l_41[4369]    = ( l_42 [4640] & !i[1820]) | ( l_42 [4641] &  i[1820]);
assign l_41[4370]    = ( l_42 [4642] & !i[1820]) | ( l_42 [4643] &  i[1820]);
assign l_41[4371]    = ( l_42 [4644] & !i[1820]) | ( l_42 [4645] &  i[1820]);
assign l_41[4372]    = ( l_42 [4646] & !i[1820]) | ( l_42 [4647] &  i[1820]);
assign l_41[4373]    = ( l_42 [4648] & !i[1820]) | ( l_42 [4649] &  i[1820]);
assign l_41[4374]    = ( l_42 [4650] & !i[1820]) | ( l_42 [4651] &  i[1820]);
assign l_41[4375]    = ( l_42 [4652] & !i[1820]) | ( l_42 [4653] &  i[1820]);
assign l_41[4376]    = ( l_42 [4654] & !i[1820]) | ( l_42 [4655] &  i[1820]);
assign l_41[4377]    = ( l_42 [4656] & !i[1820]) | ( l_42 [4657] &  i[1820]);
assign l_41[4378]    = ( l_42 [4658] & !i[1820]) | ( l_42 [4659] &  i[1820]);
assign l_41[4379]    = ( l_42 [4660] & !i[1820]) | ( l_42 [4661] &  i[1820]);
assign l_41[4380]    = ( l_42 [4662] & !i[1820]) | ( l_42 [4663] &  i[1820]);
assign l_41[4381]    = ( l_42 [4664] & !i[1820]) | ( l_42 [4665] &  i[1820]);
assign l_41[4382]    = ( l_42 [4666] & !i[1820]) | ( l_42 [4667] &  i[1820]);
assign l_41[4383]    = ( l_42 [4668] & !i[1820]) | ( l_42 [4669] &  i[1820]);
assign l_41[4384]    = ( l_42 [4670] & !i[1820]) | ( l_42 [4671] &  i[1820]);
assign l_41[4385]    = ( l_42 [4672] & !i[1820]) | ( l_42 [4673] &  i[1820]);
assign l_41[4386]    = ( l_42 [4674] & !i[1820]) | ( l_42 [4675] &  i[1820]);
assign l_41[4387]    = ( l_42 [4676] & !i[1820]) | ( l_42 [4677] &  i[1820]);
assign l_41[4388]    = ( l_42 [4678] & !i[1820]) | ( l_42 [4679] &  i[1820]);
assign l_41[4389]    = ( l_42 [4680] & !i[1820]) | ( l_42 [4681] &  i[1820]);
assign l_41[4390]    = ( l_42 [4682] & !i[1820]) | ( l_42 [4683] &  i[1820]);
assign l_41[4391]    = ( l_42 [4684] & !i[1820]) | ( l_42 [4685] &  i[1820]);
assign l_41[4392]    = ( l_42 [4686] & !i[1820]) | ( l_42 [4687] &  i[1820]);
assign l_41[4393]    = ( l_42 [4688] & !i[1820]) | ( l_42 [4689] &  i[1820]);
assign l_41[4394]    = ( l_42 [4690] & !i[1820]) | ( l_42 [4691] &  i[1820]);
assign l_41[4395]    = ( l_42 [4692] & !i[1820]) | ( l_42 [4693] &  i[1820]);
assign l_41[4396]    = ( l_42 [4694] & !i[1820]) | ( l_42 [4695] &  i[1820]);
assign l_41[4397]    = ( l_42 [4696] & !i[1820]) | ( l_42 [4697] &  i[1820]);
assign l_41[4398]    = ( l_42 [4698] & !i[1820]) | ( l_42 [4699] &  i[1820]);
assign l_41[4399]    = ( l_42 [4700] & !i[1820]) | ( l_42 [4701] &  i[1820]);
assign l_41[4400]    = ( l_42 [4702] & !i[1820]) | ( l_42 [4703] &  i[1820]);
assign l_41[4401]    = ( l_42 [4704] & !i[1820]) | ( l_42 [4705] &  i[1820]);
assign l_41[4402]    = ( l_42 [4706] & !i[1820]) | ( l_42 [4707] &  i[1820]);
assign l_41[4403]    = ( l_42 [4708] & !i[1820]) | ( l_42 [4709] &  i[1820]);
assign l_41[4404]    = ( l_42 [4710] & !i[1820]) | ( l_42 [4711] &  i[1820]);
assign l_41[4405]    = ( l_42 [4712] & !i[1820]) | ( l_42 [4713] &  i[1820]);
assign l_41[4406]    = ( l_42 [4714] & !i[1820]) | ( l_42 [4715] &  i[1820]);
assign l_41[4407]    = ( l_42 [4716] & !i[1820]) | ( l_42 [4717] &  i[1820]);
assign l_41[4408]    = ( l_42 [4718] & !i[1820]) | ( l_42 [4719] &  i[1820]);
assign l_41[4409]    = ( l_42 [4720] & !i[1820]) | ( l_42 [4721] &  i[1820]);
assign l_41[4410]    = ( l_42 [4722] & !i[1820]) | ( l_42 [4723] &  i[1820]);
assign l_41[4411]    = ( l_42 [4724] & !i[1820]) | ( l_42 [4725] &  i[1820]);
assign l_41[4412]    = ( l_42 [4726] & !i[1820]) | ( l_42 [4727] &  i[1820]);
assign l_41[4413]    = ( l_42 [4728] & !i[1820]) | ( l_42 [4729] &  i[1820]);
assign l_41[4414]    = ( l_42 [4730] & !i[1820]) | ( l_42 [4731] &  i[1820]);
assign l_41[4415]    = ( l_42 [4732] & !i[1820]) | ( l_42 [4733] &  i[1820]);
assign l_41[4416]    = ( l_42 [4734] & !i[1820]) | ( l_42 [4735] &  i[1820]);
assign l_41[4417]    = ( l_42 [4736] & !i[1820]) | ( l_42 [4737] &  i[1820]);
assign l_41[4418]    = ( l_42 [4738] & !i[1820]) | ( l_42 [4739] &  i[1820]);
assign l_41[4419]    = ( l_42 [4740] & !i[1820]) | ( l_42 [4741] &  i[1820]);
assign l_41[4420]    = ( l_42 [4742] & !i[1820]) | ( l_42 [4743] &  i[1820]);
assign l_41[4421]    = ( l_42 [4744] & !i[1820]) | ( l_42 [4745] &  i[1820]);
assign l_41[4422]    = ( l_42 [4746] & !i[1820]) | ( l_42 [4747] &  i[1820]);
assign l_41[4423]    = ( l_42 [4748] & !i[1820]) | ( l_42 [4749] &  i[1820]);
assign l_41[4424]    = ( l_42 [4750] & !i[1820]) | ( l_42 [4751] &  i[1820]);
assign l_41[4425]    = ( l_42 [4752] & !i[1820]) | ( l_42 [4753] &  i[1820]);
assign l_41[4426]    = ( l_42 [4754] & !i[1820]) | ( l_42 [4755] &  i[1820]);
assign l_41[4427]    = ( l_42 [4756] & !i[1820]) | ( l_42 [4757] &  i[1820]);
assign l_41[4428]    = ( l_42 [4758] & !i[1820]) | ( l_42 [4759] &  i[1820]);
assign l_41[4429]    = ( l_42 [4760] & !i[1820]) | ( l_42 [4761] &  i[1820]);
assign l_41[4430]    = ( l_42 [4762] & !i[1820]) | ( l_42 [4763] &  i[1820]);
assign l_41[4431]    = ( l_42 [4764] & !i[1820]) | ( l_42 [4765] &  i[1820]);
assign l_41[4432]    = ( l_42 [4766] & !i[1820]) | ( l_42 [4767] &  i[1820]);
assign l_41[4433]    = ( l_42 [4768] & !i[1820]) | ( l_42 [4769] &  i[1820]);
assign l_41[4434]    = ( l_42 [4770] & !i[1820]) | ( l_42 [4771] &  i[1820]);
assign l_41[4435]    = ( l_42 [4772] & !i[1820]) | ( l_42 [4773] &  i[1820]);
assign l_41[4436]    = ( l_42 [4774] & !i[1820]) | ( l_42 [4775] &  i[1820]);
assign l_41[4437]    = ( l_42 [4776] & !i[1820]) | ( l_42 [4777] &  i[1820]);
assign l_41[4438]    = ( l_42 [4778] & !i[1820]) | ( l_42 [4779] &  i[1820]);
assign l_41[4439]    = ( l_42 [4780] & !i[1820]) | ( l_42 [4781] &  i[1820]);
assign l_41[4440]    = ( l_42 [4782] & !i[1820]) | ( l_42 [4783] &  i[1820]);
assign l_41[4441]    = ( l_42 [4784] & !i[1820]) | ( l_42 [4785] &  i[1820]);
assign l_41[4442]    = ( l_42 [4786] & !i[1820]) | ( l_42 [4787] &  i[1820]);
assign l_41[4443]    = ( l_42 [4788] & !i[1820]) | ( l_42 [4789] &  i[1820]);
assign l_41[4444]    = ( l_42 [4790] & !i[1820]) | ( l_42 [4791] &  i[1820]);
assign l_41[4445]    = ( l_42 [4792] & !i[1820]) | ( l_42 [4793] &  i[1820]);
assign l_41[4446]    = ( l_42 [4794] & !i[1820]) | ( l_42 [4795] &  i[1820]);
assign l_41[4447]    = ( l_42 [4796] & !i[1820]) | ( l_42 [4797] &  i[1820]);
assign l_41[4448]    = ( l_42 [4798] & !i[1820]) | ( l_42 [4799] &  i[1820]);
assign l_41[4449]    = ( l_42 [4800] & !i[1820]) | ( l_42 [4801] &  i[1820]);
assign l_41[4450]    = ( l_42 [4802] & !i[1820]) | ( l_42 [4803] &  i[1820]);
assign l_41[4451]    = ( l_42 [4804] & !i[1820]) | ( l_42 [4805] &  i[1820]);
assign l_41[4452]    = ( l_42 [4806] & !i[1820]) | ( l_42 [4807] &  i[1820]);
assign l_41[4453]    = ( l_42 [4808] & !i[1820]) | ( l_42 [4809] &  i[1820]);
assign l_41[4454]    = ( l_42 [4810] & !i[1820]) | ( l_42 [4811] &  i[1820]);
assign l_41[4455]    = ( l_42 [4812] & !i[1820]) | ( l_42 [4813] &  i[1820]);
assign l_41[4456]    = ( l_42 [4814] & !i[1820]) | ( l_42 [4815] &  i[1820]);
assign l_41[4457]    = ( l_42 [4816] & !i[1820]) | ( l_42 [4817] &  i[1820]);
assign l_41[4458]    = ( l_42 [4818] & !i[1820]) | ( l_42 [4819] &  i[1820]);
assign l_41[4459]    = ( l_42 [4820] & !i[1820]) | ( l_42 [4821] &  i[1820]);
assign l_41[4460]    = ( l_42 [4822] & !i[1820]) | ( l_42 [4823] &  i[1820]);
assign l_41[4461]    = ( l_42 [4824] & !i[1820]) | ( l_42 [4825] &  i[1820]);
assign l_41[4462]    = ( l_42 [4826] & !i[1820]) | ( l_42 [4827] &  i[1820]);
assign l_41[4463]    = ( l_42 [4828] & !i[1820]) | ( l_42 [4829] &  i[1820]);
assign l_41[4464]    = ( l_42 [4830] & !i[1820]) | ( l_42 [4831] &  i[1820]);
assign l_41[4465]    = ( l_42 [4832] & !i[1820]) | ( l_42 [4833] &  i[1820]);
assign l_41[4466]    = ( l_42 [4834] & !i[1820]) | ( l_42 [4835] &  i[1820]);
assign l_41[4467]    = ( l_42 [4836] & !i[1820]) | ( l_42 [4837] &  i[1820]);
assign l_41[4468]    = ( l_42 [4838] & !i[1820]) | ( l_42 [4839] &  i[1820]);
assign l_41[4469]    = ( l_42 [4840] & !i[1820]) | ( l_42 [4841] &  i[1820]);
assign l_41[4470]    = ( l_42 [4842] & !i[1820]) | ( l_42 [4843] &  i[1820]);
assign l_41[4471]    = ( l_42 [4844] & !i[1820]) | ( l_42 [4845] &  i[1820]);
assign l_41[4472]    = ( l_42 [4846] & !i[1820]) | ( l_42 [4847] &  i[1820]);
assign l_41[4473]    = ( l_42 [4848] & !i[1820]) | ( l_42 [4849] &  i[1820]);
assign l_41[4474]    = ( l_42 [4850] & !i[1820]) | ( l_42 [4851] &  i[1820]);
assign l_41[4475]    = ( l_42 [4852] & !i[1820]) | ( l_42 [4853] &  i[1820]);
assign l_41[4476]    = ( l_42 [4854] & !i[1820]) | ( l_42 [4855] &  i[1820]);
assign l_41[4477]    = ( l_42 [4856] & !i[1820]) | ( l_42 [4857] &  i[1820]);
assign l_41[4478]    = ( l_42 [4858] & !i[1820]) | ( l_42 [4859] &  i[1820]);
assign l_41[4479]    = ( l_42 [4860] & !i[1820]) | ( l_42 [4861] &  i[1820]);
assign l_41[4480]    = ( l_42 [4862] & !i[1820]) | ( l_42 [4863] &  i[1820]);
assign l_41[4481]    = ( l_42 [4864] & !i[1820]) | ( l_42 [4865] &  i[1820]);
assign l_41[4482]    = ( l_42 [4866] & !i[1820]) | ( l_42 [4867] &  i[1820]);
assign l_41[4483]    = ( l_42 [4868] & !i[1820]) | ( l_42 [4869] &  i[1820]);
assign l_41[4484]    = ( l_42 [4870] & !i[1820]) | ( l_42 [4871] &  i[1820]);
assign l_41[4485]    = ( l_42 [4872] & !i[1820]) | ( l_42 [4873] &  i[1820]);
assign l_41[4486]    = ( l_42 [4874] & !i[1820]) | ( l_42 [4875] &  i[1820]);
assign l_41[4487]    = ( l_42 [4876] & !i[1820]) | ( l_42 [4877] &  i[1820]);
assign l_41[4488]    = ( l_42 [4878] & !i[1820]) | ( l_42 [4879] &  i[1820]);
assign l_41[4489]    = ( l_42 [4880] & !i[1820]) | ( l_42 [4881] &  i[1820]);
assign l_41[4490]    = ( l_42 [4882] & !i[1820]) | ( l_42 [4883] &  i[1820]);
assign l_41[4491]    = ( l_42 [4884] & !i[1820]) | ( l_42 [4885] &  i[1820]);
assign l_41[4492]    = ( l_42 [4886] & !i[1820]) | ( l_42 [4887] &  i[1820]);
assign l_41[4493]    = ( l_42 [4888] & !i[1820]) | ( l_42 [4889] &  i[1820]);
assign l_41[4494]    = ( l_42 [4890] & !i[1820]) | ( l_42 [4891] &  i[1820]);
assign l_41[4495]    = ( l_42 [4892] & !i[1820]) | ( l_42 [4893] &  i[1820]);
assign l_41[4496]    = ( l_42 [4894] & !i[1820]) | ( l_42 [4895] &  i[1820]);
assign l_41[4497]    = ( l_42 [4896] & !i[1820]) | ( l_42 [4897] &  i[1820]);
assign l_41[4498]    = ( l_42 [4898] & !i[1820]) | ( l_42 [4899] &  i[1820]);
assign l_41[4499]    = ( l_42 [4900] & !i[1820]) | ( l_42 [4901] &  i[1820]);
assign l_41[4500]    = ( l_42 [4902] & !i[1820]) | ( l_42 [4903] &  i[1820]);
assign l_41[4501]    = ( l_42 [4904] & !i[1820]) | ( l_42 [4905] &  i[1820]);
assign l_41[4502]    = ( l_42 [4906] & !i[1820]) | ( l_42 [4907] &  i[1820]);
assign l_41[4503]    = ( l_42 [4908] & !i[1820]) | ( l_42 [4909] &  i[1820]);
assign l_41[4504]    = ( l_42 [4910] & !i[1820]) | ( l_42 [4911] &  i[1820]);
assign l_41[4505]    = ( l_42 [4912] & !i[1820]) | ( l_42 [4913] &  i[1820]);
assign l_41[4506]    = ( l_42 [4914] & !i[1820]) | ( l_42 [4915] &  i[1820]);
assign l_41[4507]    = ( l_42 [4916] & !i[1820]) | ( l_42 [4917] &  i[1820]);
assign l_41[4508]    = ( l_42 [4918] & !i[1820]) | ( l_42 [4919] &  i[1820]);
assign l_41[4509]    = ( l_42 [4920] & !i[1820]) | ( l_42 [4921] &  i[1820]);
assign l_41[4510]    = ( l_42 [4922] & !i[1820]) | ( l_42 [4923] &  i[1820]);
assign l_41[4511]    = ( l_42 [4924] & !i[1820]) | ( l_42 [4925] &  i[1820]);
assign l_41[4512]    = ( l_42 [4926] & !i[1820]) | ( l_42 [4927] &  i[1820]);
assign l_41[4513]    = ( l_42 [4928] & !i[1820]) | ( l_42 [4929] &  i[1820]);
assign l_41[4514]    = ( l_42 [4930] & !i[1820]) | ( l_42 [4931] &  i[1820]);
assign l_41[4515]    = ( l_42 [4932] & !i[1820]) | ( l_42 [4933] &  i[1820]);
assign l_41[4516]    = ( l_42 [4934] & !i[1820]) | ( l_42 [4935] &  i[1820]);
assign l_41[4517]    = ( l_42 [4936] & !i[1820]) | ( l_42 [4937] &  i[1820]);
assign l_41[4518]    = ( l_42 [4938] & !i[1820]) | ( l_42 [4939] &  i[1820]);
assign l_41[4519]    = ( l_42 [4940] & !i[1820]) | ( l_42 [4941] &  i[1820]);
assign l_41[4520]    = ( l_42 [4942] & !i[1820]) | ( l_42 [4943] &  i[1820]);
assign l_41[4521]    = ( l_42 [4944] & !i[1820]) | ( l_42 [4945] &  i[1820]);
assign l_41[4522]    = ( l_42 [4946] & !i[1820]) | ( l_42 [4947] &  i[1820]);
assign l_41[4523]    = ( l_42 [4948] & !i[1820]) | ( l_42 [4949] &  i[1820]);
assign l_41[4524]    = ( l_42 [4950] & !i[1820]) | ( l_42 [4951] &  i[1820]);
assign l_41[4525]    = ( l_42 [4952] & !i[1820]) | ( l_42 [4953] &  i[1820]);
assign l_41[4526]    = ( l_42 [4954] & !i[1820]) | ( l_42 [4955] &  i[1820]);
assign l_41[4527]    = ( l_42 [4956] & !i[1820]) | ( l_42 [4957] &  i[1820]);
assign l_41[4528]    = ( l_42 [4958] & !i[1820]) | ( l_42 [4959] &  i[1820]);
assign l_41[4529]    = ( l_42 [4960] & !i[1820]) | ( l_42 [4961] &  i[1820]);
assign l_41[4530]    = ( l_42 [4962] & !i[1820]) | ( l_42 [4963] &  i[1820]);
assign l_41[4531]    = ( l_42 [4964] & !i[1820]) | ( l_42 [4965] &  i[1820]);
assign l_41[4532]    = ( l_42 [4966] & !i[1820]) | ( l_42 [4967] &  i[1820]);
assign l_41[4533]    = ( l_42 [4968] & !i[1820]) | ( l_42 [4969] &  i[1820]);
assign l_41[4534]    = ( l_42 [4970] & !i[1820]) | ( l_42 [4971] &  i[1820]);
assign l_41[4535]    = ( l_42 [4972] & !i[1820]) | ( l_42 [4973] &  i[1820]);
assign l_41[4536]    = ( l_42 [4974] & !i[1820]) | ( l_42 [4975] &  i[1820]);
assign l_41[4537]    = ( l_42 [4976] & !i[1820]) | ( l_42 [4977] &  i[1820]);
assign l_41[4538]    = ( l_42 [4978] & !i[1820]) | ( l_42 [4979] &  i[1820]);
assign l_41[4539]    = ( l_42 [4980] & !i[1820]) | ( l_42 [4981] &  i[1820]);
assign l_41[4540]    = ( l_42 [4982] & !i[1820]) | ( l_42 [4983] &  i[1820]);
assign l_41[4541]    = ( l_42 [4984] & !i[1820]) | ( l_42 [4985] &  i[1820]);
assign l_41[4542]    = ( l_42 [4986] & !i[1820]) | ( l_42 [4987] &  i[1820]);
assign l_41[4543]    = ( l_42 [4988] & !i[1820]) | ( l_42 [4989] &  i[1820]);
assign l_41[4544]    = ( l_42 [4990] & !i[1820]) | ( l_42 [4991] &  i[1820]);
assign l_41[4545]    = ( l_42 [4992] & !i[1820]) | ( l_42 [4993] &  i[1820]);
assign l_41[4546]    = ( l_42 [4994] & !i[1820]) | ( l_42 [4995] &  i[1820]);
assign l_41[4547]    = ( l_42 [4996] & !i[1820]) | ( l_42 [4997] &  i[1820]);
assign l_41[4548]    = ( l_42 [4998] & !i[1820]) | ( l_42 [4999] &  i[1820]);
assign l_41[4549]    = ( l_42 [5000] & !i[1820]) | ( l_42 [5001] &  i[1820]);
assign l_41[4550]    = ( l_42 [5002] & !i[1820]) | ( l_42 [5003] &  i[1820]);
assign l_41[4551]    = ( l_42 [5004] & !i[1820]) | ( l_42 [5005] &  i[1820]);
assign l_41[4552]    = ( l_42 [5006] & !i[1820]) | ( l_42 [5007] &  i[1820]);
assign l_41[4553]    = ( l_42 [5008] & !i[1820]) | ( l_42 [5009] &  i[1820]);
assign l_41[4554]    = ( l_42 [5010] & !i[1820]) | ( l_42 [5011] &  i[1820]);
assign l_41[4555]    = ( l_42 [5012] & !i[1820]) | ( l_42 [5013] &  i[1820]);
assign l_41[4556]    = ( l_42 [5014] & !i[1820]) | ( l_42 [5015] &  i[1820]);
assign l_41[4557]    = ( l_42 [5016] & !i[1820]) | ( l_42 [5017] &  i[1820]);
assign l_41[4558]    = ( l_42 [5018] & !i[1820]) | ( l_42 [5019] &  i[1820]);
assign l_41[4559]    = ( l_42 [5020] & !i[1820]) | ( l_42 [5021] &  i[1820]);
assign l_41[4560]    = ( l_42 [5022] & !i[1820]) | ( l_42 [5023] &  i[1820]);
assign l_41[4561]    = ( l_42 [5024] & !i[1820]) | ( l_42 [5025] &  i[1820]);
assign l_41[4562]    = ( l_42 [5026] & !i[1820]) | ( l_42 [5027] &  i[1820]);
assign l_41[4563]    = ( l_42 [5028] & !i[1820]) | ( l_42 [5029] &  i[1820]);
assign l_41[4564]    = ( l_42 [5030] & !i[1820]) | ( l_42 [5031] &  i[1820]);
assign l_41[4565]    = ( l_42 [5032] & !i[1820]) | ( l_42 [5033] &  i[1820]);
assign l_41[4566]    = ( l_42 [5034] & !i[1820]) | ( l_42 [5035] &  i[1820]);
assign l_41[4567]    = ( l_42 [5036] & !i[1820]) | ( l_42 [5037] &  i[1820]);
assign l_41[4568]    = ( l_42 [5038] & !i[1820]) | ( l_42 [5039] &  i[1820]);
assign l_41[4569]    = ( l_42 [5040] & !i[1820]) | ( l_42 [5041] &  i[1820]);
assign l_41[4570]    = ( l_42 [5042] & !i[1820]) | ( l_42 [5043] &  i[1820]);
assign l_41[4571]    = ( l_42 [5044] & !i[1820]) | ( l_42 [5045] &  i[1820]);
assign l_41[4572]    = ( l_42 [5046] & !i[1820]) | ( l_42 [5047] &  i[1820]);
assign l_41[4573]    = ( l_42 [5048] & !i[1820]) | ( l_42 [5049] &  i[1820]);
assign l_41[4574]    = ( l_42 [5050] & !i[1820]) | ( l_42 [5051] &  i[1820]);
assign l_41[4575]    = ( l_42 [5052] & !i[1820]) | ( l_42 [5053] &  i[1820]);
assign l_41[4576]    = ( l_42 [5054] & !i[1820]) | ( l_42 [5055] &  i[1820]);
assign l_41[4577]    = ( l_42 [5056] & !i[1820]) | ( l_42 [5057] &  i[1820]);
assign l_41[4578]    = ( l_42 [5058] & !i[1820]) | ( l_42 [5059] &  i[1820]);
assign l_41[4579]    = ( l_42 [5060] & !i[1820]) | ( l_42 [5061] &  i[1820]);
assign l_41[4580]    = ( l_42 [5062] & !i[1820]) | ( l_42 [5063] &  i[1820]);
assign l_41[4581]    = ( l_42 [5064] & !i[1820]) | ( l_42 [5065] &  i[1820]);
assign l_41[4582]    = ( l_42 [5066] & !i[1820]) | ( l_42 [5067] &  i[1820]);
assign l_41[4583]    = ( l_42 [5068] & !i[1820]) | ( l_42 [5069] &  i[1820]);
assign l_41[4584]    = ( l_42 [5070] & !i[1820]) | ( l_42 [5071] &  i[1820]);
assign l_41[4585]    = ( l_42 [5072] & !i[1820]) | ( l_42 [5073] &  i[1820]);
assign l_41[4586]    = ( l_42 [5074] & !i[1820]) | ( l_42 [5075] &  i[1820]);
assign l_41[4587]    = ( l_42 [5076] & !i[1820]) | ( l_42 [5077] &  i[1820]);
assign l_41[4588]    = ( l_42 [5078] & !i[1820]) | ( l_42 [5079] &  i[1820]);
assign l_41[4589]    = ( l_42 [5080] & !i[1820]) | ( l_42 [5081] &  i[1820]);
assign l_41[4590]    = ( l_42 [5082] & !i[1820]) | ( l_42 [5083] &  i[1820]);
assign l_41[4591]    = ( l_42 [5084] & !i[1820]) | ( l_42 [5085] &  i[1820]);
assign l_41[4592]    = ( l_42 [5086] & !i[1820]) | ( l_42 [5087] &  i[1820]);
assign l_41[4593]    = ( l_42 [5088] & !i[1820]) | ( l_42 [5089] &  i[1820]);
assign l_41[4594]    = ( l_42 [5090] & !i[1820]) | ( l_42 [5091] &  i[1820]);
assign l_41[4595]    = ( l_42 [5092] & !i[1820]) | ( l_42 [5093] &  i[1820]);
assign l_41[4596]    = ( l_42 [5094] & !i[1820]) | ( l_42 [5095] &  i[1820]);
assign l_41[4597]    = ( l_42 [5096] & !i[1820]) | ( l_42 [5097] &  i[1820]);
assign l_41[4598]    = ( l_42 [5098] & !i[1820]) | ( l_42 [5099] &  i[1820]);
assign l_41[4599]    = ( l_42 [5100] & !i[1820]) | ( l_42 [5101] &  i[1820]);
assign l_41[4600]    = ( l_42 [5102] & !i[1820]) | ( l_42 [5103] &  i[1820]);
assign l_41[4601]    = ( l_42 [5104] & !i[1820]) | ( l_42 [5105] &  i[1820]);
assign l_41[4602]    = ( l_42 [5106] & !i[1820]) | ( l_42 [5107] &  i[1820]);
assign l_41[4603]    = ( l_42 [5108] & !i[1820]) | ( l_42 [5109] &  i[1820]);
assign l_41[4604]    = ( l_42 [5110] & !i[1820]) | ( l_42 [5111] &  i[1820]);
assign l_41[4605]    = ( l_42 [5112] & !i[1820]) | ( l_42 [5113] &  i[1820]);
assign l_41[4606]    = ( l_42 [5114] & !i[1820]) | ( l_42 [5115] &  i[1820]);
assign l_41[4607]    = ( l_42 [5116] & !i[1820]) | ( l_42 [5117] &  i[1820]);
assign l_41[4608]    = ( l_42 [5118] & !i[1820]) | ( l_42 [5119] &  i[1820]);
assign l_41[4609]    = ( l_42 [5120] & !i[1820]) | ( l_42 [5121] &  i[1820]);
assign l_41[4610]    = ( l_42 [5122] & !i[1820]) | ( l_42 [5123] &  i[1820]);
assign l_41[4611]    = ( l_42 [5124] & !i[1820]) | ( l_42 [5125] &  i[1820]);
assign l_41[4612]    = ( l_42 [5126] & !i[1820]) | ( l_42 [5127] &  i[1820]);
assign l_41[4613]    = ( l_42 [5128] & !i[1820]) | ( l_42 [5129] &  i[1820]);
assign l_41[4614]    = ( l_42 [5130] & !i[1820]) | ( l_42 [5131] &  i[1820]);
assign l_41[4615]    = ( l_42 [5132] & !i[1820]) | ( l_42 [5133] &  i[1820]);
assign l_41[4616]    = ( l_42 [5134] & !i[1820]) | ( l_42 [5135] &  i[1820]);
assign l_41[4617]    = ( l_42 [5136] & !i[1820]) | ( l_42 [5137] &  i[1820]);
assign l_41[4618]    = ( l_42 [5138] & !i[1820]) | ( l_42 [5139] &  i[1820]);
assign l_41[4619]    = ( l_42 [5140] & !i[1820]) | ( l_42 [5141] &  i[1820]);
assign l_41[4620]    = ( l_42 [5142] & !i[1820]) | ( l_42 [5143] &  i[1820]);
assign l_41[4621]    = ( l_42 [5144] & !i[1820]) | ( l_42 [5145] &  i[1820]);
assign l_41[4622]    = ( l_42 [5146] & !i[1820]) | ( l_42 [5147] &  i[1820]);
assign l_41[4623]    = ( l_42 [5148] & !i[1820]) | ( l_42 [5149] &  i[1820]);
assign l_41[4624]    = ( l_42 [5150] & !i[1820]) | ( l_42 [5151] &  i[1820]);
assign l_41[4625]    = ( l_42 [5152] & !i[1820]) | ( l_42 [5153] &  i[1820]);
assign l_41[4626]    = ( l_42 [5154] & !i[1820]) | ( l_42 [5155] &  i[1820]);
assign l_41[4627]    = ( l_42 [5156] & !i[1820]) | ( l_42 [5157] &  i[1820]);
assign l_41[4628]    = ( l_42 [5158] & !i[1820]) | ( l_42 [5159] &  i[1820]);
assign l_41[4629]    = ( l_42 [5160] & !i[1820]) | ( l_42 [5161] &  i[1820]);
assign l_41[4630]    = ( l_42 [5162] & !i[1820]) | ( l_42 [5163] &  i[1820]);
assign l_41[4631]    = ( l_42 [5164] & !i[1820]) | ( l_42 [5165] &  i[1820]);
assign l_41[4632]    = ( l_42 [5166] & !i[1820]) | ( l_42 [5167] &  i[1820]);
assign l_41[4633]    = ( l_42 [5168] & !i[1820]) | ( l_42 [5169] &  i[1820]);
assign l_41[4634]    = ( l_42 [5170] & !i[1820]) | ( l_42 [5171] &  i[1820]);
assign l_41[4635]    = ( l_42 [5172] & !i[1820]) | ( l_42 [5173] &  i[1820]);
assign l_41[4636]    = ( l_42 [5174] & !i[1820]) | ( l_42 [5175] &  i[1820]);
assign l_41[4637]    = ( l_42 [5176] & !i[1820]) | ( l_42 [5177] &  i[1820]);
assign l_41[4638]    = ( l_42 [5178] & !i[1820]) | ( l_42 [5179] &  i[1820]);
assign l_41[4639]    = ( l_42 [5180] & !i[1820]) | ( l_42 [5181] &  i[1820]);
assign l_41[4640]    = ( l_42 [5182] & !i[1820]) | ( l_42 [5183] &  i[1820]);
assign l_41[4641]    = ( l_42 [5184] & !i[1820]) | ( l_42 [5185] &  i[1820]);
assign l_41[4642]    = ( l_42 [5186] & !i[1820]) | ( l_42 [5187] &  i[1820]);
assign l_41[4643]    = ( l_42 [5188] & !i[1820]) | ( l_42 [5189] &  i[1820]);
assign l_41[4644]    = ( l_42 [5190] & !i[1820]) | ( l_42 [5191] &  i[1820]);
assign l_41[4645]    = ( l_42 [5192] & !i[1820]) | ( l_42 [5193] &  i[1820]);
assign l_41[4646]    = ( l_42 [5194] & !i[1820]) | ( l_42 [5195] &  i[1820]);
assign l_41[4647]    = ( l_42 [5196] & !i[1820]) | ( l_42 [5197] &  i[1820]);
assign l_41[4648]    = ( l_42 [5198] & !i[1820]) | ( l_42 [5199] &  i[1820]);
assign l_41[4649]    = ( l_42 [5200] & !i[1820]) | ( l_42 [5201] &  i[1820]);
assign l_41[4650]    = ( l_42 [5202] & !i[1820]) | ( l_42 [5203] &  i[1820]);
assign l_41[4651]    = ( l_42 [5204] & !i[1820]) | ( l_42 [5205] &  i[1820]);
assign l_41[4652]    = ( l_42 [5206] & !i[1820]) | ( l_42 [5207] &  i[1820]);
assign l_41[4653]    = ( l_42 [5208] & !i[1820]) | ( l_42 [5209] &  i[1820]);
assign l_41[4654]    = ( l_42 [5210] & !i[1820]) | ( l_42 [5211] &  i[1820]);
assign l_41[4655]    = ( l_42 [5212] & !i[1820]) | ( l_42 [5213] &  i[1820]);
assign l_41[4656]    = ( l_42 [5214] & !i[1820]) | ( l_42 [5215] &  i[1820]);
assign l_41[4657]    = ( l_42 [5216] & !i[1820]) | ( l_42 [5217] &  i[1820]);
assign l_41[4658]    = ( l_42 [5218] & !i[1820]) | ( l_42 [5219] &  i[1820]);
assign l_41[4659]    = ( l_42 [5220] & !i[1820]) | ( l_42 [5221] &  i[1820]);
assign l_41[4660]    = ( l_42 [5222] & !i[1820]) | ( l_42 [5223] &  i[1820]);
assign l_41[4661]    = ( l_42 [5224] & !i[1820]) | ( l_42 [5225] &  i[1820]);
assign l_41[4662]    = ( l_42 [5226] & !i[1820]) | ( l_42 [5227] &  i[1820]);
assign l_41[4663]    = ( l_42 [5228] & !i[1820]) | ( l_42 [5229] &  i[1820]);
assign l_41[4664]    = ( l_42 [5230] & !i[1820]) | ( l_42 [5231] &  i[1820]);
assign l_41[4665]    = ( l_42 [5232] & !i[1820]) | ( l_42 [5233] &  i[1820]);
assign l_41[4666]    = ( l_42 [5234] & !i[1820]) | ( l_42 [5235] &  i[1820]);
assign l_41[4667]    = ( l_42 [5236] & !i[1820]) | ( l_42 [5237] &  i[1820]);
assign l_41[4668]    = ( l_42 [5238] & !i[1820]) | ( l_42 [5239] &  i[1820]);
assign l_41[4669]    = ( l_42 [5240] & !i[1820]) | ( l_42 [5241] &  i[1820]);
assign l_41[4670]    = ( l_42 [5242] & !i[1820]) | ( l_42 [5243] &  i[1820]);
assign l_41[4671]    = ( l_42 [5244] & !i[1820]) | ( l_42 [5245] &  i[1820]);
assign l_41[4672]    = ( l_42 [5246] & !i[1820]) | ( l_42 [5247] &  i[1820]);
assign l_41[4673]    = ( l_42 [5248] & !i[1820]) | ( l_42 [5249] &  i[1820]);
assign l_41[4674]    = ( l_42 [5250] & !i[1820]) | ( l_42 [5251] &  i[1820]);
assign l_41[4675]    = ( l_42 [5252] & !i[1820]) | ( l_42 [5253] &  i[1820]);
assign l_41[4676]    = ( l_42 [5254] & !i[1820]) | ( l_42 [5255] &  i[1820]);
assign l_41[4677]    = ( l_42 [5256] & !i[1820]) | ( l_42 [5257] &  i[1820]);
assign l_41[4678]    = ( l_42 [5258] & !i[1820]) | ( l_42 [5259] &  i[1820]);
assign l_41[4679]    = ( l_42 [5260] & !i[1820]) | ( l_42 [5261] &  i[1820]);
assign l_41[4680]    = ( l_42 [5262] & !i[1820]) | ( l_42 [5263] &  i[1820]);
assign l_41[4681]    = ( l_42 [5264] & !i[1820]) | ( l_42 [5265] &  i[1820]);
assign l_41[4682]    = ( l_42 [5266] & !i[1820]) | ( l_42 [5267] &  i[1820]);
assign l_41[4683]    = ( l_42 [5268] & !i[1820]) | ( l_42 [5269] &  i[1820]);
assign l_41[4684]    = ( l_42 [5270] & !i[1820]) | ( l_42 [5271] &  i[1820]);
assign l_41[4685]    = ( l_42 [5272] & !i[1820]) | ( l_42 [5273] &  i[1820]);
assign l_41[4686]    = ( l_42 [5274] & !i[1820]) | ( l_42 [5275] &  i[1820]);
assign l_41[4687]    = ( l_42 [5276] & !i[1820]) | ( l_42 [5277] &  i[1820]);
assign l_41[4688]    = ( l_42 [5278] & !i[1820]) | ( l_42 [5279] &  i[1820]);
assign l_41[4689]    = ( l_42 [5280] & !i[1820]) | ( l_42 [5281] &  i[1820]);
assign l_41[4690]    = ( l_42 [5282] & !i[1820]) | ( l_42 [5283] &  i[1820]);
assign l_41[4691]    = ( l_42 [5284] & !i[1820]) | ( l_42 [5285] &  i[1820]);
assign l_41[4692]    = ( l_42 [5286] & !i[1820]) | ( l_42 [5287] &  i[1820]);
assign l_41[4693]    = ( l_42 [5288] & !i[1820]) | ( l_42 [5289] &  i[1820]);
assign l_41[4694]    = ( l_42 [5290] & !i[1820]) | ( l_42 [5291] &  i[1820]);
assign l_41[4695]    = ( l_42 [5292] & !i[1820]) | ( l_42 [5293] &  i[1820]);
assign l_41[4696]    = ( l_42 [5294] & !i[1820]) | ( l_42 [5295] &  i[1820]);
assign l_41[4697]    = ( l_42 [5296] & !i[1820]) | ( l_42 [5297] &  i[1820]);
assign l_41[4698]    = ( l_42 [5298] & !i[1820]) | ( l_42 [5299] &  i[1820]);
assign l_41[4699]    = ( l_42 [5300] & !i[1820]) | ( l_42 [5301] &  i[1820]);
assign l_41[4700]    = ( l_42 [5302] & !i[1820]) | ( l_42 [5303] &  i[1820]);
assign l_41[4701]    = ( l_42 [5304] & !i[1820]) | ( l_42 [5305] &  i[1820]);
assign l_41[4702]    = ( l_42 [5306] & !i[1820]) | ( l_42 [5307] &  i[1820]);
assign l_41[4703]    = ( l_42 [5308] & !i[1820]) | ( l_42 [5309] &  i[1820]);
assign l_41[4704]    = ( l_42 [5310] & !i[1820]) | ( l_42 [5311] &  i[1820]);
assign l_41[4705]    = ( l_42 [5312] & !i[1820]) | ( l_42 [5313] &  i[1820]);
assign l_41[4706]    = ( l_42 [5314] & !i[1820]) | ( l_42 [5315] &  i[1820]);
assign l_41[4707]    = ( l_42 [5316] & !i[1820]) | ( l_42 [5317] &  i[1820]);
assign l_41[4708]    = ( l_42 [5318] & !i[1820]) | ( l_42 [5319] &  i[1820]);
assign l_41[4709]    = ( l_42 [5320] & !i[1820]) | ( l_42 [5321] &  i[1820]);
assign l_41[4710]    = ( l_42 [5322] & !i[1820]) | ( l_42 [5323] &  i[1820]);
assign l_41[4711]    = ( l_42 [5324] & !i[1820]) | ( l_42 [5325] &  i[1820]);
assign l_41[4712]    = ( l_42 [5326] & !i[1820]) | ( l_42 [5327] &  i[1820]);
assign l_41[4713]    = ( l_42 [5328] & !i[1820]) | ( l_42 [5329] &  i[1820]);
assign l_41[4714]    = ( l_42 [5330] & !i[1820]) | ( l_42 [5331] &  i[1820]);
assign l_41[4715]    = ( l_42 [5332] & !i[1820]) | ( l_42 [5333] &  i[1820]);
assign l_41[4716]    = ( l_42 [5334] & !i[1820]) | ( l_42 [5335] &  i[1820]);
assign l_41[4717]    = ( l_42 [5336] & !i[1820]) | ( l_42 [5337] &  i[1820]);
assign l_41[4718]    = ( l_42 [5338] & !i[1820]) | ( l_42 [5339] &  i[1820]);
assign l_41[4719]    = ( l_42 [5340] & !i[1820]) | ( l_42 [5341] &  i[1820]);
assign l_41[4720]    = ( l_42 [5342] & !i[1820]) | ( l_42 [5343] &  i[1820]);
assign l_41[4721]    = ( l_42 [5344] & !i[1820]) | ( l_42 [5345] &  i[1820]);
assign l_41[4722]    = ( l_42 [5346] & !i[1820]) | ( l_42 [5347] &  i[1820]);
assign l_41[4723]    = ( l_42 [5348] & !i[1820]) | ( l_42 [5349] &  i[1820]);
assign l_41[4724]    = ( l_42 [5350] & !i[1820]) | ( l_42 [5351] &  i[1820]);
assign l_41[4725]    = ( l_42 [5352] & !i[1820]) | ( l_42 [5353] &  i[1820]);
assign l_41[4726]    = ( l_42 [5354] & !i[1820]) | ( l_42 [5355] &  i[1820]);
assign l_41[4727]    = ( l_42 [5356] & !i[1820]) | ( l_42 [5357] &  i[1820]);
assign l_41[4728]    = ( l_42 [5358] & !i[1820]) | ( l_42 [5359] &  i[1820]);
assign l_41[4729]    = ( l_42 [5360] & !i[1820]) | ( l_42 [5361] &  i[1820]);
assign l_41[4730]    = ( l_42 [5362] & !i[1820]) | ( l_42 [5363] &  i[1820]);
assign l_41[4731]    = ( l_42 [5364] & !i[1820]) | ( l_42 [5365] &  i[1820]);
assign l_41[4732]    = ( l_42 [5366] & !i[1820]) | ( l_42 [5367] &  i[1820]);
assign l_41[4733]    = ( l_42 [5368] & !i[1820]) | ( l_42 [5369] &  i[1820]);
assign l_41[4734]    = ( l_42 [5370] & !i[1820]) | ( l_42 [5371] &  i[1820]);
assign l_41[4735]    = ( l_42 [5372] & !i[1820]) | ( l_42 [5373] &  i[1820]);
assign l_41[4736]    = ( l_42 [5374] & !i[1820]) | ( l_42 [5375] &  i[1820]);
assign l_41[4737]    = ( l_42 [5376] & !i[1820]) | ( l_42 [5377] &  i[1820]);
assign l_41[4738]    = ( l_42 [5378] & !i[1820]) | ( l_42 [5379] &  i[1820]);
assign l_41[4739]    = ( l_42 [5380] & !i[1820]) | ( l_42 [5381] &  i[1820]);
assign l_41[4740]    = ( l_42 [5382] & !i[1820]) | ( l_42 [5383] &  i[1820]);
assign l_41[4741]    = ( l_42 [5384] & !i[1820]) | ( l_42 [5385] &  i[1820]);
assign l_41[4742]    = ( l_42 [5386] & !i[1820]) | ( l_42 [5387] &  i[1820]);
assign l_41[4743]    = ( l_42 [5388] & !i[1820]) | ( l_42 [5389] &  i[1820]);
assign l_41[4744]    = ( l_42 [5390] & !i[1820]) | ( l_42 [5391] &  i[1820]);
assign l_41[4745]    = ( l_42 [5392] & !i[1820]) | ( l_42 [5393] &  i[1820]);
assign l_41[4746]    = ( l_42 [5394] & !i[1820]) | ( l_42 [5395] &  i[1820]);
assign l_41[4747]    = ( l_42 [5396] & !i[1820]) | ( l_42 [5397] &  i[1820]);
assign l_41[4748]    = ( l_42 [5398] & !i[1820]) | ( l_42 [5399] &  i[1820]);
assign l_41[4749]    = ( l_42 [5400] & !i[1820]) | ( l_42 [5401] &  i[1820]);
assign l_41[4750]    = ( l_42 [5402] & !i[1820]) | ( l_42 [5403] &  i[1820]);
assign l_41[4751]    = ( l_42 [5404] & !i[1820]) | ( l_42 [5405] &  i[1820]);
assign l_41[4752]    = ( l_42 [5406] & !i[1820]) | ( l_42 [5407] &  i[1820]);
assign l_41[4753]    = ( l_42 [5408] & !i[1820]) | ( l_42 [5409] &  i[1820]);
assign l_41[4754]    = ( l_42 [5410] & !i[1820]) | ( l_42 [5411] &  i[1820]);
assign l_41[4755]    = ( l_42 [5412] & !i[1820]) | ( l_42 [5413] &  i[1820]);
assign l_41[4756]    = ( l_42 [5414] & !i[1820]) | ( l_42 [5415] &  i[1820]);
assign l_41[4757]    = ( l_42 [5416] & !i[1820]) | ( l_42 [5417] &  i[1820]);
assign l_41[4758]    = ( l_42 [5418] & !i[1820]) | ( l_42 [5419] &  i[1820]);
assign l_41[4759]    = ( l_42 [5420] & !i[1820]) | ( l_42 [5421] &  i[1820]);
assign l_41[4760]    = ( l_42 [5422] & !i[1820]) | ( l_42 [5423] &  i[1820]);
assign l_41[4761]    = ( l_42 [5424] & !i[1820]) | ( l_42 [5425] &  i[1820]);
assign l_41[4762]    = ( l_42 [5426] & !i[1820]) | ( l_42 [5427] &  i[1820]);
assign l_41[4763]    = ( l_42 [5428] & !i[1820]) | ( l_42 [5429] &  i[1820]);
assign l_41[4764]    = ( l_42 [5430] & !i[1820]) | ( l_42 [5431] &  i[1820]);
assign l_41[4765]    = ( l_42 [5432] & !i[1820]) | ( l_42 [5433] &  i[1820]);
assign l_41[4766]    = ( l_42 [5434] & !i[1820]) | ( l_42 [5435] &  i[1820]);
assign l_41[4767]    = ( l_42 [5436] & !i[1820]) | ( l_42 [5437] &  i[1820]);
assign l_41[4768]    = ( l_42 [5438] & !i[1820]) | ( l_42 [5439] &  i[1820]);
assign l_41[4769]    = ( l_42 [5440] & !i[1820]) | ( l_42 [5441] &  i[1820]);
assign l_41[4770]    = ( l_42 [5442] & !i[1820]) | ( l_42 [5443] &  i[1820]);
assign l_41[4771]    = ( l_42 [5444] & !i[1820]) | ( l_42 [5445] &  i[1820]);
assign l_41[4772]    = ( l_42 [5446] & !i[1820]) | ( l_42 [5447] &  i[1820]);
assign l_41[4773]    = ( l_42 [5448] & !i[1820]) | ( l_42 [5449] &  i[1820]);
assign l_41[4774]    = ( l_42 [5450] & !i[1820]) | ( l_42 [5451] &  i[1820]);
assign l_41[4775]    = ( l_42 [5452] & !i[1820]) | ( l_42 [5453] &  i[1820]);
assign l_41[4776]    = ( l_42 [5454] & !i[1820]) | ( l_42 [5455] &  i[1820]);
assign l_41[4777]    = ( l_42 [5456] & !i[1820]) | ( l_42 [5457] &  i[1820]);
assign l_41[4778]    = ( l_42 [5458] & !i[1820]) | ( l_42 [5459] &  i[1820]);
assign l_41[4779]    = ( l_42 [5460] & !i[1820]) | ( l_42 [5461] &  i[1820]);
assign l_41[4780]    = ( l_42 [5462] & !i[1820]) | ( l_42 [5463] &  i[1820]);
assign l_41[4781]    = ( l_42 [5464] & !i[1820]) | ( l_42 [5465] &  i[1820]);
assign l_41[4782]    = ( l_42 [5466] & !i[1820]) | ( l_42 [5467] &  i[1820]);
assign l_41[4783]    = ( l_42 [5468] & !i[1820]) | ( l_42 [5469] &  i[1820]);
assign l_41[4784]    = ( l_42 [5470] & !i[1820]) | ( l_42 [5471] &  i[1820]);
assign l_41[4785]    = ( l_42 [5472] & !i[1820]) | ( l_42 [5473] &  i[1820]);
assign l_41[4786]    = ( l_42 [5474] & !i[1820]) | ( l_42 [5475] &  i[1820]);
assign l_41[4787]    = ( l_42 [5476] & !i[1820]) | ( l_42 [5477] &  i[1820]);
assign l_41[4788]    = ( l_42 [5478] & !i[1820]) | ( l_42 [5479] &  i[1820]);
assign l_41[4789]    = ( l_42 [5480] & !i[1820]) | ( l_42 [5481] &  i[1820]);
assign l_41[4790]    = ( l_42 [5482] & !i[1820]) | ( l_42 [5483] &  i[1820]);
assign l_41[4791]    = ( l_42 [5484] & !i[1820]) | ( l_42 [5485] &  i[1820]);
assign l_41[4792]    = ( l_42 [5486] & !i[1820]) | ( l_42 [5487] &  i[1820]);
assign l_41[4793]    = ( l_42 [5488] & !i[1820]) | ( l_42 [5489] &  i[1820]);
assign l_41[4794]    = ( l_42 [5490] & !i[1820]) | ( l_42 [5491] &  i[1820]);
assign l_41[4795]    = ( l_42 [5492] & !i[1820]) | ( l_42 [5493] &  i[1820]);
assign l_41[4796]    = ( l_42 [5494] & !i[1820]) | ( l_42 [5495] &  i[1820]);
assign l_41[4797]    = ( l_42 [5496] & !i[1820]) | ( l_42 [5497] &  i[1820]);
assign l_41[4798]    = ( l_42 [5498] & !i[1820]) | ( l_42 [5499] &  i[1820]);
assign l_41[4799]    = ( l_42 [5500] & !i[1820]) | ( l_42 [5501] &  i[1820]);
assign l_41[4800]    = ( l_42 [5502] & !i[1820]) | ( l_42 [5503] &  i[1820]);
assign l_41[4801]    = ( l_42 [5504] & !i[1820]) | ( l_42 [5505] &  i[1820]);
assign l_41[4802]    = ( l_42 [5506] & !i[1820]) | ( l_42 [5507] &  i[1820]);
assign l_41[4803]    = ( l_42 [5508] & !i[1820]) | ( l_42 [5509] &  i[1820]);
assign l_41[4804]    = ( l_42 [5510] & !i[1820]) | ( l_42 [5511] &  i[1820]);
assign l_41[4805]    = ( l_42 [5512] & !i[1820]) | ( l_42 [5513] &  i[1820]);
assign l_41[4806]    = ( l_42 [5514] & !i[1820]) | ( l_42 [5515] &  i[1820]);
assign l_41[4807]    = ( l_42 [5516] & !i[1820]) | ( l_42 [5517] &  i[1820]);
assign l_41[4808]    = ( l_42 [5518] & !i[1820]) | ( l_42 [5519] &  i[1820]);
assign l_41[4809]    = ( l_42 [5520] & !i[1820]) | ( l_42 [5521] &  i[1820]);
assign l_41[4810]    = ( l_42 [5522] & !i[1820]) | ( l_42 [5523] &  i[1820]);
assign l_41[4811]    = ( l_42 [5524] & !i[1820]) | ( l_42 [5525] &  i[1820]);
assign l_41[4812]    = ( l_42 [5526] & !i[1820]) | ( l_42 [5527] &  i[1820]);
assign l_41[4813]    = ( l_42 [5528] & !i[1820]) | ( l_42 [5529] &  i[1820]);
assign l_41[4814]    = ( l_42 [5530] & !i[1820]) | ( l_42 [5531] &  i[1820]);
assign l_41[4815]    = ( l_42 [5532] & !i[1820]) | ( l_42 [5533] &  i[1820]);
assign l_41[4816]    = ( l_42 [5534] & !i[1820]) | ( l_42 [5535] &  i[1820]);
assign l_41[4817]    = ( l_42 [5536] & !i[1820]) | ( l_42 [5537] &  i[1820]);
assign l_41[4818]    = ( l_42 [5538] & !i[1820]) | ( l_42 [5539] &  i[1820]);
assign l_41[4819]    = ( l_42 [5540] & !i[1820]) | ( l_42 [5541] &  i[1820]);
assign l_41[4820]    = ( l_42 [5542] & !i[1820]) | ( l_42 [5543] &  i[1820]);
assign l_41[4821]    = ( l_42 [5544] & !i[1820]) | ( l_42 [5545] &  i[1820]);
assign l_41[4822]    = ( l_42 [5546] & !i[1820]) | ( l_42 [5547] &  i[1820]);
assign l_41[4823]    = ( l_42 [5548] & !i[1820]) | ( l_42 [5549] &  i[1820]);
assign l_41[4824]    = ( l_42 [5550] & !i[1820]) | ( l_42 [5551] &  i[1820]);
assign l_41[4825]    = ( l_42 [5552] & !i[1820]) | ( l_42 [5553] &  i[1820]);
assign l_41[4826]    = ( l_42 [5554] & !i[1820]) | ( l_42 [5555] &  i[1820]);
assign l_41[4827]    = ( l_42 [5556] & !i[1820]) | ( l_42 [5557] &  i[1820]);
assign l_41[4828]    = ( l_42 [5558] & !i[1820]) | ( l_42 [5559] &  i[1820]);
assign l_41[4829]    = ( l_42 [5560] & !i[1820]) | ( l_42 [5561] &  i[1820]);
assign l_41[4830]    = ( l_42 [5562] & !i[1820]) | ( l_42 [5563] &  i[1820]);
assign l_41[4831]    = ( l_42 [5564] & !i[1820]) | ( l_42 [5565] &  i[1820]);
assign l_41[4832]    = ( l_42 [5566] & !i[1820]) | ( l_42 [5567] &  i[1820]);
assign l_41[4833]    = ( l_42 [5568] & !i[1820]) | ( l_42 [5569] &  i[1820]);
assign l_41[4834]    = ( l_42 [5570] & !i[1820]) | ( l_42 [5571] &  i[1820]);
assign l_41[4835]    = ( l_42 [5572] & !i[1820]) | ( l_42 [5573] &  i[1820]);
assign l_41[4836]    = ( l_42 [5574] & !i[1820]) | ( l_42 [5575] &  i[1820]);
assign l_41[4837]    = ( l_42 [5576] & !i[1820]) | ( l_42 [5577] &  i[1820]);
assign l_41[4838]    = ( l_42 [5578] & !i[1820]) | ( l_42 [5579] &  i[1820]);
assign l_41[4839]    = ( l_42 [5580] & !i[1820]) | ( l_42 [5581] &  i[1820]);
assign l_41[4840]    = ( l_42 [5582] & !i[1820]) | ( l_42 [5583] &  i[1820]);
assign l_41[4841]    = ( l_42 [5584] & !i[1820]) | ( l_42 [5585] &  i[1820]);
assign l_41[4842]    = ( l_42 [5586] & !i[1820]) | ( l_42 [5587] &  i[1820]);
assign l_41[4843]    = ( l_42 [5588] & !i[1820]) | ( l_42 [5589] &  i[1820]);
assign l_41[4844]    = ( l_42 [5590] & !i[1820]) | ( l_42 [5591] &  i[1820]);
assign l_41[4845]    = ( l_42 [5592] & !i[1820]) | ( l_42 [5593] &  i[1820]);
assign l_41[4846]    = ( l_42 [5594] & !i[1820]) | ( l_42 [5595] &  i[1820]);
assign l_41[4847]    = ( l_42 [5596] & !i[1820]) | ( l_42 [5597] &  i[1820]);
assign l_41[4848]    = ( l_42 [5598] & !i[1820]) | ( l_42 [5599] &  i[1820]);
assign l_41[4849]    = ( l_42 [5600] & !i[1820]) | ( l_42 [5601] &  i[1820]);
assign l_41[4850]    = ( l_42 [5602] & !i[1820]) | ( l_42 [5603] &  i[1820]);
assign l_41[4851]    = ( l_42 [5604] & !i[1820]) | ( l_42 [5605] &  i[1820]);
assign l_41[4852]    = ( l_42 [5606] & !i[1820]) | ( l_42 [5607] &  i[1820]);
assign l_41[4853]    = ( l_42 [5608] & !i[1820]) | ( l_42 [5609] &  i[1820]);
assign l_41[4854]    = ( l_42 [5610] & !i[1820]) | ( l_42 [5611] &  i[1820]);
assign l_41[4855]    = ( l_42 [5612] & !i[1820]) | ( l_42 [5613] &  i[1820]);
assign l_41[4856]    = ( l_42 [5614] & !i[1820]) | ( l_42 [5615] &  i[1820]);
assign l_41[4857]    = ( l_42 [5616] & !i[1820]) | ( l_42 [5617] &  i[1820]);
assign l_41[4858]    = ( l_42 [5618] & !i[1820]) | ( l_42 [5619] &  i[1820]);
assign l_41[4859]    = ( l_42 [5620] & !i[1820]) | ( l_42 [5621] &  i[1820]);
assign l_41[4860]    = ( l_42 [5622] & !i[1820]) | ( l_42 [5623] &  i[1820]);
assign l_41[4861]    = ( l_42 [5624] & !i[1820]) | ( l_42 [5625] &  i[1820]);
assign l_41[4862]    = ( l_42 [5626] & !i[1820]) | ( l_42 [5627] &  i[1820]);
assign l_41[4863]    = ( l_42 [5628] & !i[1820]) | ( l_42 [5629] &  i[1820]);
assign l_41[4864]    = ( l_42 [5630] & !i[1820]) | ( l_42 [5631] &  i[1820]);
assign l_41[4865]    = ( l_42 [5632] & !i[1820]) | ( l_42 [5633] &  i[1820]);
assign l_41[4866]    = ( l_42 [5634] & !i[1820]) | ( l_42 [5635] &  i[1820]);
assign l_41[4867]    = ( l_42 [5636] & !i[1820]) | ( l_42 [5637] &  i[1820]);
assign l_41[4868]    = ( l_42 [5638] & !i[1820]) | ( l_42 [5639] &  i[1820]);
assign l_41[4869]    = ( l_42 [5640] & !i[1820]) | ( l_42 [5641] &  i[1820]);
assign l_41[4870]    = ( l_42 [5642] & !i[1820]) | ( l_42 [5643] &  i[1820]);
assign l_41[4871]    = ( l_42 [5644] & !i[1820]) | ( l_42 [5645] &  i[1820]);
assign l_41[4872]    = ( l_42 [5646] & !i[1820]) | ( l_42 [5647] &  i[1820]);
assign l_41[4873]    = ( l_42 [5648] & !i[1820]) | ( l_42 [5649] &  i[1820]);
assign l_41[4874]    = ( l_42 [5650] & !i[1820]) | ( l_42 [5651] &  i[1820]);
assign l_41[4875]    = ( l_42 [5652] & !i[1820]) | ( l_42 [5653] &  i[1820]);
assign l_41[4876]    = ( l_42 [5654] & !i[1820]) | ( l_42 [5655] &  i[1820]);
assign l_41[4877]    = ( l_42 [5656] & !i[1820]) | ( l_42 [5657] &  i[1820]);
assign l_41[4878]    = ( l_42 [5658] & !i[1820]) | ( l_42 [5659] &  i[1820]);
assign l_41[4879]    = ( l_42 [5660] & !i[1820]) | ( l_42 [5661] &  i[1820]);
assign l_41[4880]    = ( l_42 [5662] & !i[1820]) | ( l_42 [5663] &  i[1820]);
assign l_41[4881]    = ( l_42 [5664] & !i[1820]) | ( l_42 [5665] &  i[1820]);
assign l_41[4882]    = ( l_42 [5666] & !i[1820]) | ( l_42 [5667] &  i[1820]);
assign l_41[4883]    = ( l_42 [5668] & !i[1820]) | ( l_42 [5669] &  i[1820]);
assign l_41[4884]    = ( l_42 [5670] & !i[1820]) | ( l_42 [5671] &  i[1820]);
assign l_41[4885]    = ( l_42 [5672] & !i[1820]) | ( l_42 [5673] &  i[1820]);
assign l_41[4886]    = ( l_42 [5674] & !i[1820]) | ( l_42 [5675] &  i[1820]);
assign l_41[4887]    = ( l_42 [5676] & !i[1820]) | ( l_42 [5677] &  i[1820]);
assign l_41[4888]    = ( l_42 [5678] & !i[1820]) | ( l_42 [5679] &  i[1820]);
assign l_41[4889]    = ( l_42 [5680] & !i[1820]) | ( l_42 [5681] &  i[1820]);
assign l_41[4890]    = ( l_42 [5682] & !i[1820]) | ( l_42 [5683] &  i[1820]);
assign l_41[4891]    = ( l_42 [5684] & !i[1820]) | ( l_42 [5685] &  i[1820]);
assign l_41[4892]    = ( l_42 [5686] & !i[1820]) | ( l_42 [5687] &  i[1820]);
assign l_41[4893]    = ( l_42 [5688] & !i[1820]) | ( l_42 [5689] &  i[1820]);
assign l_41[4894]    = ( l_42 [5690] & !i[1820]) | ( l_42 [5691] &  i[1820]);
assign l_41[4895]    = ( l_42 [5692] & !i[1820]) | ( l_42 [5693] &  i[1820]);
assign l_41[4896]    = ( l_42 [5694] & !i[1820]) | ( l_42 [5695] &  i[1820]);
assign l_41[4897]    = ( l_42 [5696] & !i[1820]) | ( l_42 [5697] &  i[1820]);
assign l_41[4898]    = ( l_42 [5698] & !i[1820]) | ( l_42 [5699] &  i[1820]);
assign l_41[4899]    = ( l_42 [5700] & !i[1820]) | ( l_42 [5701] &  i[1820]);
assign l_41[4900]    = ( l_42 [5702] & !i[1820]) | ( l_42 [5703] &  i[1820]);
assign l_41[4901]    = ( l_42 [5704] & !i[1820]) | ( l_42 [5705] &  i[1820]);
assign l_41[4902]    = ( l_42 [5706] & !i[1820]) | ( l_42 [5707] &  i[1820]);
assign l_41[4903]    = ( l_42 [5708] & !i[1820]) | ( l_42 [5709] &  i[1820]);
assign l_41[4904]    = ( l_42 [5710] & !i[1820]) | ( l_42 [5711] &  i[1820]);
assign l_41[4905]    = ( l_42 [5712] & !i[1820]) | ( l_42 [5713] &  i[1820]);
assign l_41[4906]    = ( l_42 [5714] & !i[1820]) | ( l_42 [5715] &  i[1820]);
assign l_41[4907]    = ( l_42 [5716] & !i[1820]) | ( l_42 [5717] &  i[1820]);
assign l_41[4908]    = ( l_42 [5718] & !i[1820]) | ( l_42 [5719] &  i[1820]);
assign l_41[4909]    = ( l_42 [5720] & !i[1820]) | ( l_42 [5721] &  i[1820]);
assign l_41[4910]    = ( l_42 [5722] & !i[1820]) | ( l_42 [5723] &  i[1820]);
assign l_41[4911]    = ( l_42 [5724] & !i[1820]) | ( l_42 [5725] &  i[1820]);
assign l_41[4912]    = ( l_42 [5726] & !i[1820]) | ( l_42 [5727] &  i[1820]);
assign l_41[4913]    = ( l_42 [5728] & !i[1820]) | ( l_42 [5729] &  i[1820]);
assign l_41[4914]    = ( l_42 [5730] & !i[1820]) | ( l_42 [5731] &  i[1820]);
assign l_41[4915]    = ( l_42 [5732] & !i[1820]) | ( l_42 [5733] &  i[1820]);
assign l_41[4916]    = ( l_42 [5734] & !i[1820]) | ( l_42 [5735] &  i[1820]);
assign l_41[4917]    = ( l_42 [5736] & !i[1820]) | ( l_42 [5737] &  i[1820]);
assign l_41[4918]    = ( l_42 [5738] & !i[1820]) | ( l_42 [5739] &  i[1820]);
assign l_41[4919]    = ( l_42 [5740] & !i[1820]) | ( l_42 [5741] &  i[1820]);
assign l_41[4920]    = ( l_42 [5742] & !i[1820]) | ( l_42 [5743] &  i[1820]);
assign l_41[4921]    = ( l_42 [5744] & !i[1820]) | ( l_42 [5745] &  i[1820]);
assign l_41[4922]    = ( l_42 [5746] & !i[1820]) | ( l_42 [5747] &  i[1820]);
assign l_41[4923]    = ( l_42 [5748] & !i[1820]) | ( l_42 [5749] &  i[1820]);
assign l_41[4924]    = ( l_42 [5750] & !i[1820]) | ( l_42 [5751] &  i[1820]);
assign l_41[4925]    = ( l_42 [5752] & !i[1820]) | ( l_42 [5753] &  i[1820]);
assign l_41[4926]    = ( l_42 [5754] & !i[1820]) | ( l_42 [5755] &  i[1820]);
assign l_41[4927]    = ( l_42 [5756] & !i[1820]) | ( l_42 [5757] &  i[1820]);
assign l_41[4928]    = ( l_42 [5758] & !i[1820]) | ( l_42 [5759] &  i[1820]);
assign l_41[4929]    = ( l_42 [5760] & !i[1820]) | ( l_42 [5761] &  i[1820]);
assign l_41[4930]    = ( l_42 [5762] & !i[1820]) | ( l_42 [5763] &  i[1820]);
assign l_41[4931]    = ( l_42 [5764] & !i[1820]) | ( l_42 [5765] &  i[1820]);
assign l_41[4932]    = ( l_42 [5766] & !i[1820]) | ( l_42 [5767] &  i[1820]);
assign l_41[4933]    = ( l_42 [5768] & !i[1820]) | ( l_42 [5769] &  i[1820]);
assign l_41[4934]    = ( l_42 [5770] & !i[1820]) | ( l_42 [5771] &  i[1820]);
assign l_41[4935]    = ( l_42 [5772] & !i[1820]) | ( l_42 [5773] &  i[1820]);
assign l_41[4936]    = ( l_42 [5774] & !i[1820]) | ( l_42 [5775] &  i[1820]);
assign l_41[4937]    = ( l_42 [5776] & !i[1820]) | ( l_42 [5777] &  i[1820]);
assign l_41[4938]    = ( l_42 [5778] & !i[1820]) | ( l_42 [5779] &  i[1820]);
assign l_41[4939]    = ( l_42 [5780] & !i[1820]) | ( l_42 [5781] &  i[1820]);
assign l_41[4940]    = ( l_42 [5782] & !i[1820]) | ( l_42 [5783] &  i[1820]);
assign l_41[4941]    = ( l_42 [5784] & !i[1820]) | ( l_42 [5785] &  i[1820]);
assign l_41[4942]    = ( l_42 [5786] & !i[1820]) | ( l_42 [5787] &  i[1820]);
assign l_41[4943]    = ( l_42 [5788] & !i[1820]) | ( l_42 [5789] &  i[1820]);
assign l_41[4944]    = ( l_42 [5790] & !i[1820]) | ( l_42 [5791] &  i[1820]);
assign l_41[4945]    = ( l_42 [5792] & !i[1820]) | ( l_42 [5793] &  i[1820]);
assign l_41[4946]    = ( l_42 [5794] & !i[1820]) | ( l_42 [5795] &  i[1820]);
assign l_41[4947]    = ( l_42 [5796] & !i[1820]) | ( l_42 [5797] &  i[1820]);
assign l_41[4948]    = ( l_42 [5798] & !i[1820]) | ( l_42 [5799] &  i[1820]);
assign l_41[4949]    = ( l_42 [5800] & !i[1820]) | ( l_42 [5801] &  i[1820]);
assign l_41[4950]    = ( l_42 [5802] & !i[1820]) | ( l_42 [5803] &  i[1820]);
assign l_41[4951]    = ( l_42 [5804] & !i[1820]) | ( l_42 [5805] &  i[1820]);
assign l_41[4952]    = ( l_42 [5806] & !i[1820]) | ( l_42 [5807] &  i[1820]);
assign l_41[4953]    = ( l_42 [5808] & !i[1820]) | ( l_42 [5809] &  i[1820]);
assign l_41[4954]    = ( l_42 [5810] & !i[1820]) | ( l_42 [5811] &  i[1820]);
assign l_41[4955]    = ( l_42 [5812] & !i[1820]) | ( l_42 [5813] &  i[1820]);
assign l_41[4956]    = ( l_42 [5814] & !i[1820]) | ( l_42 [5815] &  i[1820]);
assign l_41[4957]    = ( l_42 [5816] & !i[1820]) | ( l_42 [5817] &  i[1820]);
assign l_41[4958]    = ( l_42 [5818] & !i[1820]) | ( l_42 [5819] &  i[1820]);
assign l_41[4959]    = ( l_42 [5820] & !i[1820]) | ( l_42 [5821] &  i[1820]);
assign l_41[4960]    = ( l_42 [5822] & !i[1820]) | ( l_42 [5823] &  i[1820]);
assign l_41[4961]    = ( l_42 [5824] & !i[1820]) | ( l_42 [5825] &  i[1820]);
assign l_41[4962]    = ( l_42 [5826] & !i[1820]) | ( l_42 [5827] &  i[1820]);
assign l_41[4963]    = ( l_42 [5828] & !i[1820]) | ( l_42 [5829] &  i[1820]);
assign l_41[4964]    = ( l_42 [5830] & !i[1820]) | ( l_42 [5831] &  i[1820]);
assign l_41[4965]    = ( l_42 [5832] & !i[1820]) | ( l_42 [5833] &  i[1820]);
assign l_41[4966]    = ( l_42 [5834] & !i[1820]) | ( l_42 [5835] &  i[1820]);
assign l_41[4967]    = ( l_42 [5836] & !i[1820]) | ( l_42 [5837] &  i[1820]);
assign l_41[4968]    = ( l_42 [5838] & !i[1820]) | ( l_42 [5839] &  i[1820]);
assign l_41[4969]    = ( l_42 [5840] & !i[1820]) | ( l_42 [5841] &  i[1820]);
assign l_41[4970]    = ( l_42 [5842] & !i[1820]) | ( l_42 [5843] &  i[1820]);
assign l_41[4971]    = ( l_42 [5844] & !i[1820]) | ( l_42 [5845] &  i[1820]);
assign l_41[4972]    = ( l_42 [5846] & !i[1820]) | ( l_42 [5847] &  i[1820]);
assign l_41[4973]    = ( l_42 [5848] & !i[1820]) | ( l_42 [5849] &  i[1820]);
assign l_41[4974]    = ( l_42 [5850] & !i[1820]) | ( l_42 [5851] &  i[1820]);
assign l_41[4975]    = ( l_42 [5852] & !i[1820]) | ( l_42 [5853] &  i[1820]);
assign l_41[4976]    = ( l_42 [5854] & !i[1820]) | ( l_42 [5855] &  i[1820]);
assign l_41[4977]    = ( l_42 [5856] & !i[1820]) | ( l_42 [5857] &  i[1820]);
assign l_41[4978]    = ( l_42 [5858] & !i[1820]) | ( l_42 [5859] &  i[1820]);
assign l_41[4979]    = ( l_42 [5860] & !i[1820]) | ( l_42 [5861] &  i[1820]);
assign l_41[4980]    = ( l_42 [5862] & !i[1820]) | ( l_42 [5863] &  i[1820]);
assign l_41[4981]    = ( l_42 [5864] & !i[1820]) | ( l_42 [5865] &  i[1820]);
assign l_41[4982]    = ( l_42 [5866] & !i[1820]) | ( l_42 [5867] &  i[1820]);
assign l_41[4983]    = ( l_42 [5868] & !i[1820]) | ( l_42 [5869] &  i[1820]);
assign l_41[4984]    = ( l_42 [5870] & !i[1820]) | ( l_42 [5871] &  i[1820]);
assign l_41[4985]    = ( l_42 [5872] & !i[1820]) | ( l_42 [5873] &  i[1820]);
assign l_41[4986]    = ( l_42 [5874] & !i[1820]) | ( l_42 [5875] &  i[1820]);
assign l_41[4987]    = ( l_42 [5876] & !i[1820]) | ( l_42 [5877] &  i[1820]);
assign l_41[4988]    = ( l_42 [5878] & !i[1820]) | ( l_42 [5879] &  i[1820]);
assign l_41[4989]    = ( l_42 [5880] & !i[1820]) | ( l_42 [5881] &  i[1820]);
assign l_41[4990]    = ( l_42 [5882] & !i[1820]) | ( l_42 [5883] &  i[1820]);
assign l_41[4991]    = ( l_42 [5884] & !i[1820]) | ( l_42 [5885] &  i[1820]);
assign l_41[4992]    = ( l_42 [5886] & !i[1820]) | ( l_42 [5887] &  i[1820]);
assign l_41[4993]    = ( l_42 [5888] & !i[1820]) | ( l_42 [5889] &  i[1820]);
assign l_41[4994]    = ( l_42 [5890] & !i[1820]) | ( l_42 [5891] &  i[1820]);
assign l_41[4995]    = ( l_42 [5892] & !i[1820]) | ( l_42 [5893] &  i[1820]);
assign l_41[4996]    = ( l_42 [5894] & !i[1820]) | ( l_42 [5895] &  i[1820]);
assign l_41[4997]    = ( l_42 [5896] & !i[1820]) | ( l_42 [5897] &  i[1820]);
assign l_41[4998]    = ( l_42 [5898] & !i[1820]) | ( l_42 [5899] &  i[1820]);
assign l_41[4999]    = ( l_42 [5900] & !i[1820]) | ( l_42 [5901] &  i[1820]);
assign l_41[5000]    = ( l_42 [5902] & !i[1820]) | ( l_42 [5903] &  i[1820]);
assign l_41[5001]    = ( l_42 [5904] & !i[1820]) | ( l_42 [5905] &  i[1820]);
assign l_41[5002]    = ( l_42 [5906] & !i[1820]) | ( l_42 [5907] &  i[1820]);
assign l_41[5003]    = ( l_42 [5908] & !i[1820]) | ( l_42 [5909] &  i[1820]);
assign l_41[5004]    = ( l_42 [5910] & !i[1820]) | ( l_42 [5911] &  i[1820]);
assign l_41[5005]    = ( l_42 [5912] & !i[1820]) | ( l_42 [5913] &  i[1820]);
assign l_41[5006]    = ( l_42 [5914] & !i[1820]) | ( l_42 [5915] &  i[1820]);
assign l_41[5007]    = ( l_42 [5916] & !i[1820]) | ( l_42 [5917] &  i[1820]);
assign l_41[5008]    = ( l_42 [5918] & !i[1820]) | ( l_42 [5919] &  i[1820]);
assign l_41[5009]    = ( l_42 [5920] & !i[1820]) | ( l_42 [5921] &  i[1820]);
assign l_41[5010]    = ( l_42 [5922] & !i[1820]) | ( l_42 [5923] &  i[1820]);
assign l_41[5011]    = ( l_42 [5924] & !i[1820]) | ( l_42 [5925] &  i[1820]);
assign l_41[5012]    = ( l_42 [5926] & !i[1820]) | ( l_42 [5927] &  i[1820]);
assign l_41[5013]    = ( l_42 [5928] & !i[1820]) | ( l_42 [5929] &  i[1820]);
assign l_41[5014]    = ( l_42 [5930] & !i[1820]) | ( l_42 [5931] &  i[1820]);
assign l_41[5015]    = ( l_42 [5932] & !i[1820]) | ( l_42 [5933] &  i[1820]);
assign l_41[5016]    = ( l_42 [5934] & !i[1820]) | ( l_42 [5935] &  i[1820]);
assign l_41[5017]    = ( l_42 [5936] & !i[1820]) | ( l_42 [5937] &  i[1820]);
assign l_41[5018]    = ( l_42 [5938] & !i[1820]) | ( l_42 [5939] &  i[1820]);
assign l_41[5019]    = ( l_42 [5940] & !i[1820]) | ( l_42 [5941] &  i[1820]);
assign l_41[5020]    = ( l_42 [5942] & !i[1820]) | ( l_42 [5943] &  i[1820]);
assign l_41[5021]    = ( l_42 [5944] & !i[1820]) | ( l_42 [5945] &  i[1820]);
assign l_41[5022]    = ( l_42 [5946] & !i[1820]) | ( l_42 [5947] &  i[1820]);
assign l_41[5023]    = ( l_42 [5948] & !i[1820]) | ( l_42 [5949] &  i[1820]);
assign l_41[5024]    = ( l_42 [5950] & !i[1820]) | ( l_42 [5951] &  i[1820]);
assign l_41[5025]    = ( l_42 [5952] & !i[1820]) | ( l_42 [5953] &  i[1820]);
assign l_41[5026]    = ( l_42 [5954] & !i[1820]) | ( l_42 [5955] &  i[1820]);
assign l_41[5027]    = ( l_42 [5956] & !i[1820]) | ( l_42 [5957] &  i[1820]);
assign l_41[5028]    = ( l_42 [5958] & !i[1820]) | ( l_42 [5959] &  i[1820]);
assign l_41[5029]    = ( l_42 [5960] & !i[1820]) | ( l_42 [5961] &  i[1820]);
assign l_41[5030]    = ( l_42 [5962] & !i[1820]) | ( l_42 [5963] &  i[1820]);
assign l_41[5031]    = ( l_42 [5964] & !i[1820]) | ( l_42 [5965] &  i[1820]);
assign l_41[5032]    = ( l_42 [5966] & !i[1820]) | ( l_42 [5967] &  i[1820]);
assign l_41[5033]    = ( l_42 [5968] & !i[1820]) | ( l_42 [5969] &  i[1820]);
assign l_41[5034]    = ( l_42 [5970] & !i[1820]) | ( l_42 [5971] &  i[1820]);
assign l_41[5035]    = ( l_42 [5972] & !i[1820]) | ( l_42 [5973] &  i[1820]);
assign l_41[5036]    = ( l_42 [5974] & !i[1820]) | ( l_42 [5975] &  i[1820]);
assign l_41[5037]    = ( l_42 [5976] & !i[1820]) | ( l_42 [5977] &  i[1820]);
assign l_41[5038]    = ( l_42 [5978] & !i[1820]) | ( l_42 [5979] &  i[1820]);
assign l_41[5039]    = ( l_42 [5980] & !i[1820]) | ( l_42 [5981] &  i[1820]);
assign l_41[5040]    = ( l_42 [5982] & !i[1820]) | ( l_42 [5983] &  i[1820]);
assign l_41[5041]    = ( l_42 [5984] & !i[1820]) | ( l_42 [5985] &  i[1820]);
assign l_41[5042]    = ( l_42 [5986] & !i[1820]) | ( l_42 [5987] &  i[1820]);
assign l_41[5043]    = ( l_42 [5988] & !i[1820]) | ( l_42 [5989] &  i[1820]);
assign l_41[5044]    = ( l_42 [5990] & !i[1820]) | ( l_42 [5991] &  i[1820]);
assign l_41[5045]    = ( l_42 [5992] & !i[1820]) | ( l_42 [5993] &  i[1820]);
assign l_41[5046]    = ( l_42 [5994] & !i[1820]) | ( l_42 [5995] &  i[1820]);
assign l_41[5047]    = ( l_42 [5996] & !i[1820]) | ( l_42 [5997] &  i[1820]);
assign l_41[5048]    = ( l_42 [5998] & !i[1820]) | ( l_42 [5999] &  i[1820]);
assign l_41[5049]    = ( l_42 [6000] & !i[1820]) | ( l_42 [6001] &  i[1820]);
assign l_41[5050]    = ( l_42 [6002] & !i[1820]) | ( l_42 [6003] &  i[1820]);
assign l_41[5051]    = ( l_42 [6004] & !i[1820]) | ( l_42 [6005] &  i[1820]);
assign l_41[5052]    = ( l_42 [6006] & !i[1820]) | ( l_42 [6007] &  i[1820]);
assign l_41[5053]    = ( l_42 [6008] & !i[1820]) | ( l_42 [6009] &  i[1820]);
assign l_41[5054]    = ( l_42 [6010] & !i[1820]) | ( l_42 [6011] &  i[1820]);
assign l_41[5055]    = ( l_42 [6012] & !i[1820]) | ( l_42 [6013] &  i[1820]);
assign l_41[5056]    = ( l_42 [6014] & !i[1820]) | ( l_42 [6015] &  i[1820]);
assign l_41[5057]    = ( l_42 [6016] & !i[1820]) | ( l_42 [6017] &  i[1820]);
assign l_41[5058]    = ( l_42 [6018] & !i[1820]) | ( l_42 [6019] &  i[1820]);
assign l_41[5059]    = ( l_42 [6020] & !i[1820]) | ( l_42 [6021] &  i[1820]);
assign l_41[5060]    = ( l_42 [6022] & !i[1820]) | ( l_42 [6023] &  i[1820]);
assign l_41[5061]    = ( l_42 [6024] & !i[1820]) | ( l_42 [6025] &  i[1820]);
assign l_41[5062]    = ( l_42 [6026] & !i[1820]) | ( l_42 [6027] &  i[1820]);
assign l_41[5063]    = ( l_42 [6028] & !i[1820]) | ( l_42 [6029] &  i[1820]);
assign l_41[5064]    = ( l_42 [6030] & !i[1820]) | ( l_42 [6031] &  i[1820]);
assign l_41[5065]    = ( l_42 [6032] & !i[1820]) | ( l_42 [6033] &  i[1820]);
assign l_41[5066]    = ( l_42 [6034] & !i[1820]) | ( l_42 [6035] &  i[1820]);
assign l_41[5067]    = ( l_42 [6036] & !i[1820]) | ( l_42 [6037] &  i[1820]);
assign l_41[5068]    = ( l_42 [6038] & !i[1820]) | ( l_42 [6039] &  i[1820]);
assign l_41[5069]    = ( l_42 [6040] & !i[1820]) | ( l_42 [6041] &  i[1820]);
assign l_41[5070]    = ( l_42 [6042] & !i[1820]) | ( l_42 [6043] &  i[1820]);
assign l_41[5071]    = ( l_42 [6044] & !i[1820]) | ( l_42 [6045] &  i[1820]);
assign l_41[5072]    = ( l_42 [6046] & !i[1820]) | ( l_42 [6047] &  i[1820]);
assign l_41[5073]    = ( l_42 [6048] & !i[1820]) | ( l_42 [6049] &  i[1820]);
assign l_41[5074]    = ( l_42 [6050] & !i[1820]) | ( l_42 [6051] &  i[1820]);
assign l_41[5075]    = ( l_42 [6052] & !i[1820]) | ( l_42 [6053] &  i[1820]);
assign l_41[5076]    = ( l_42 [6054] & !i[1820]) | ( l_42 [6055] &  i[1820]);
assign l_41[5077]    = ( l_42 [6056] & !i[1820]) | ( l_42 [6057] &  i[1820]);
assign l_41[5078]    = ( l_42 [6058] & !i[1820]) | ( l_42 [6059] &  i[1820]);
assign l_41[5079]    = ( l_42 [6060] & !i[1820]) | ( l_42 [6061] &  i[1820]);
assign l_41[5080]    = ( l_42 [6062] & !i[1820]) | ( l_42 [6063] &  i[1820]);
assign l_41[5081]    = ( l_42 [6064] & !i[1820]) | ( l_42 [6065] &  i[1820]);
assign l_41[5082]    = ( l_42 [6066] & !i[1820]) | ( l_42 [6067] &  i[1820]);
assign l_41[5083]    = ( l_42 [6068] & !i[1820]) | ( l_42 [6069] &  i[1820]);
assign l_41[5084]    = ( l_42 [6070] & !i[1820]) | ( l_42 [6071] &  i[1820]);
assign l_41[5085]    = ( l_42 [6072] & !i[1820]) | ( l_42 [6073] &  i[1820]);
assign l_41[5086]    = ( l_42 [6074] & !i[1820]) | ( l_42 [6075] &  i[1820]);
assign l_41[5087]    = ( l_42 [6076] & !i[1820]) | ( l_42 [6077] &  i[1820]);
assign l_41[5088]    = ( l_42 [6078] & !i[1820]) | ( l_42 [6079] &  i[1820]);
assign l_41[5089]    = ( l_42 [6080] & !i[1820]) | ( l_42 [6081] &  i[1820]);
assign l_41[5090]    = ( l_42 [6082] & !i[1820]) | ( l_42 [6083] &  i[1820]);
assign l_41[5091]    = ( l_42 [6084] & !i[1820]) | ( l_42 [6085] &  i[1820]);
assign l_41[5092]    = ( l_42 [6086] & !i[1820]) | ( l_42 [6087] &  i[1820]);
assign l_41[5093]    = ( l_42 [6088] & !i[1820]) | ( l_42 [6089] &  i[1820]);
assign l_41[5094]    = ( l_42 [6090] & !i[1820]) | ( l_42 [6091] &  i[1820]);
assign l_41[5095]    = ( l_42 [6092] & !i[1820]) | ( l_42 [6093] &  i[1820]);
assign l_41[5096]    = ( l_42 [6094] & !i[1820]) | ( l_42 [6095] &  i[1820]);
assign l_41[5097]    = ( l_42 [6096] & !i[1820]) | ( l_42 [6097] &  i[1820]);
assign l_41[5098]    = ( l_42 [6098] & !i[1820]) | ( l_42 [6099] &  i[1820]);
assign l_41[5099]    = ( l_42 [6100] & !i[1820]) | ( l_42 [6101] &  i[1820]);
assign l_41[5100]    = ( l_42 [6102] & !i[1820]) | ( l_42 [6103] &  i[1820]);
assign l_41[5101]    = ( l_42 [6104] & !i[1820]) | ( l_42 [6105] &  i[1820]);
assign l_41[5102]    = ( l_42 [6106] & !i[1820]) | ( l_42 [6107] &  i[1820]);
assign l_41[5103]    = ( l_42 [6108] & !i[1820]) | ( l_42 [6109] &  i[1820]);
assign l_41[5104]    = ( l_42 [6110] & !i[1820]) | ( l_42 [6111] &  i[1820]);
assign l_41[5105]    = ( l_42 [6112] & !i[1820]) | ( l_42 [6113] &  i[1820]);
assign l_41[5106]    = ( l_42 [6114] & !i[1820]) | ( l_42 [6115] &  i[1820]);
assign l_41[5107]    = ( l_42 [6116] & !i[1820]) | ( l_42 [6117] &  i[1820]);
assign l_41[5108]    = ( l_42 [6118] & !i[1820]) | ( l_42 [6119] &  i[1820]);
assign l_41[5109]    = ( l_42 [6120] & !i[1820]) | ( l_42 [6121] &  i[1820]);
assign l_41[5110]    = ( l_42 [6122] & !i[1820]) | ( l_42 [6123] &  i[1820]);
assign l_41[5111]    = ( l_42 [6124] & !i[1820]) | ( l_42 [6125] &  i[1820]);
assign l_41[5112]    = ( l_42 [6126] & !i[1820]) | ( l_42 [6127] &  i[1820]);
assign l_41[5113]    = ( l_42 [6128] & !i[1820]) | ( l_42 [6129] &  i[1820]);
assign l_41[5114]    = ( l_42 [6130] & !i[1820]) | ( l_42 [6131] &  i[1820]);
assign l_41[5115]    = ( l_42 [6132] & !i[1820]) | ( l_42 [6133] &  i[1820]);
assign l_41[5116]    = ( l_42 [6134] & !i[1820]) | ( l_42 [6135] &  i[1820]);
assign l_41[5117]    = ( l_42 [6136] & !i[1820]) | ( l_42 [6137] &  i[1820]);
assign l_41[5118]    = ( l_42 [6138] & !i[1820]) | ( l_42 [6139] &  i[1820]);
assign l_41[5119]    = ( l_42 [6140] & !i[1820]) | ( l_42 [6141] &  i[1820]);
assign l_41[5120]    = ( l_42 [6142] & !i[1820]) | ( l_42 [6143] &  i[1820]);
assign l_41[5121]    = ( l_42 [6144] & !i[1820]) | ( l_42 [6145] &  i[1820]);
assign l_41[5122]    = ( l_42 [6146] & !i[1820]) | ( l_42 [6147] &  i[1820]);
assign l_41[5123]    = ( l_42 [6148] & !i[1820]) | ( l_42 [6149] &  i[1820]);
assign l_41[5124]    = ( l_42 [6150] & !i[1820]) | ( l_42 [6151] &  i[1820]);
assign l_41[5125]    = ( l_42 [6152] & !i[1820]) | ( l_42 [6153] &  i[1820]);
assign l_41[5126]    = ( l_42 [6154] & !i[1820]) | ( l_42 [6155] &  i[1820]);
assign l_41[5127]    = ( l_42 [6156] & !i[1820]) | ( l_42 [6157] &  i[1820]);
assign l_41[5128]    = ( l_42 [6158] & !i[1820]) | ( l_42 [6159] &  i[1820]);
assign l_41[5129]    = ( l_42 [6160] & !i[1820]) | ( l_42 [6161] &  i[1820]);
assign l_41[5130]    = ( l_42 [6162] & !i[1820]) | ( l_42 [6163] &  i[1820]);
assign l_41[5131]    = ( l_42 [6164] & !i[1820]) | ( l_42 [6165] &  i[1820]);
assign l_41[5132]    = ( l_42 [6166] & !i[1820]) | ( l_42 [6167] &  i[1820]);
assign l_41[5133]    = ( l_42 [6168] & !i[1820]) | ( l_42 [6169] &  i[1820]);
assign l_41[5134]    = ( l_42 [6170] & !i[1820]) | ( l_42 [6171] &  i[1820]);
assign l_41[5135]    = ( l_42 [6172] & !i[1820]) | ( l_42 [6173] &  i[1820]);
assign l_41[5136]    = ( l_42 [6174] & !i[1820]) | ( l_42 [6175] &  i[1820]);
assign l_41[5137]    = ( l_42 [6176] & !i[1820]) | ( l_42 [6177] &  i[1820]);
assign l_41[5138]    = ( l_42 [6178] & !i[1820]) | ( l_42 [6179] &  i[1820]);
assign l_41[5139]    = ( l_42 [6180] & !i[1820]) | ( l_42 [6181] &  i[1820]);
assign l_41[5140]    = ( l_42 [6182] & !i[1820]) | ( l_42 [6183] &  i[1820]);
assign l_41[5141]    = ( l_42 [6184] & !i[1820]) | ( l_42 [6185] &  i[1820]);
assign l_41[5142]    = ( l_42 [6186] & !i[1820]) | ( l_42 [6187] &  i[1820]);
assign l_41[5143]    = ( l_42 [6188] & !i[1820]) | ( l_42 [6189] &  i[1820]);
assign l_41[5144]    = ( l_42 [6190] & !i[1820]) | ( l_42 [6191] &  i[1820]);
assign l_41[5145]    = ( l_42 [6192] & !i[1820]) | ( l_42 [6193] &  i[1820]);
assign l_41[5146]    = ( l_42 [6194] & !i[1820]) | ( l_42 [6195] &  i[1820]);
assign l_41[5147]    = ( l_42 [6196] & !i[1820]) | ( l_42 [6197] &  i[1820]);
assign l_41[5148]    = ( l_42 [6198] & !i[1820]) | ( l_42 [6199] &  i[1820]);
assign l_41[5149]    = ( l_42 [6200] & !i[1820]) | ( l_42 [6201] &  i[1820]);
assign l_41[5150]    = ( l_42 [6202] & !i[1820]) | ( l_42 [6203] &  i[1820]);
assign l_41[5151]    = ( l_42 [6204] & !i[1820]) | ( l_42 [6205] &  i[1820]);
assign l_41[5152]    = ( l_42 [6206] & !i[1820]) | ( l_42 [6207] &  i[1820]);
assign l_41[5153]    = ( l_42 [6208] & !i[1820]) | ( l_42 [6209] &  i[1820]);
assign l_41[5154]    = ( l_42 [6210] & !i[1820]) | ( l_42 [6211] &  i[1820]);
assign l_41[5155]    = ( l_42 [6212] & !i[1820]) | ( l_42 [6213] &  i[1820]);
assign l_41[5156]    = ( l_42 [6214] & !i[1820]) | ( l_42 [6215] &  i[1820]);
assign l_41[5157]    = ( l_42 [6216] & !i[1820]) | ( l_42 [6217] &  i[1820]);
assign l_41[5158]    = ( l_42 [6218] & !i[1820]) | ( l_42 [6219] &  i[1820]);
assign l_41[5159]    = ( l_42 [6220] & !i[1820]) | ( l_42 [6221] &  i[1820]);
assign l_41[5160]    = ( l_42 [6222] & !i[1820]) | ( l_42 [6223] &  i[1820]);
assign l_41[5161]    = ( l_42 [6224] & !i[1820]) | ( l_42 [6225] &  i[1820]);
assign l_41[5162]    = ( l_42 [6226] & !i[1820]) | ( l_42 [6227] &  i[1820]);
assign l_41[5163]    = ( l_42 [6228] & !i[1820]) | ( l_42 [6229] &  i[1820]);
assign l_41[5164]    = ( l_42 [6230] & !i[1820]) | ( l_42 [6231] &  i[1820]);
assign l_41[5165]    = ( l_42 [6232] & !i[1820]) | ( l_42 [6233] &  i[1820]);
assign l_41[5166]    = ( l_42 [6234] & !i[1820]) | ( l_42 [6235] &  i[1820]);
assign l_41[5167]    = ( l_42 [6236] & !i[1820]) | ( l_42 [6237] &  i[1820]);
assign l_41[5168]    = ( l_42 [6238] & !i[1820]) | ( l_42 [6239] &  i[1820]);
assign l_41[5169]    = ( l_42 [6240] & !i[1820]) | ( l_42 [6241] &  i[1820]);
assign l_41[5170]    = ( l_42 [6242] & !i[1820]) | ( l_42 [6243] &  i[1820]);
assign l_41[5171]    = ( l_42 [6244] & !i[1820]) | ( l_42 [6245] &  i[1820]);
assign l_41[5172]    = ( l_42 [6246] & !i[1820]) | ( l_42 [6247] &  i[1820]);
assign l_41[5173]    = ( l_42 [6248] & !i[1820]) | ( l_42 [6249] &  i[1820]);
assign l_41[5174]    = ( l_42 [6250] & !i[1820]) | ( l_42 [6251] &  i[1820]);
assign l_41[5175]    = ( l_42 [6252] & !i[1820]) | ( l_42 [6253] &  i[1820]);
assign l_41[5176]    = ( l_42 [6254] & !i[1820]) | ( l_42 [6255] &  i[1820]);
assign l_41[5177]    = ( l_42 [6256] & !i[1820]) | ( l_42 [6257] &  i[1820]);
assign l_41[5178]    = ( l_42 [6258] & !i[1820]) | ( l_42 [6259] &  i[1820]);
assign l_41[5179]    = ( l_42 [6260] & !i[1820]) | ( l_42 [6261] &  i[1820]);
assign l_41[5180]    = ( l_42 [6262] & !i[1820]) | ( l_42 [6263] &  i[1820]);
assign l_41[5181]    = ( l_42 [6264] & !i[1820]) | ( l_42 [6265] &  i[1820]);
assign l_41[5182]    = ( l_42 [6266] & !i[1820]) | ( l_42 [6267] &  i[1820]);
assign l_41[5183]    = ( l_42 [6268] & !i[1820]) | ( l_42 [6269] &  i[1820]);
assign l_41[5184]    = ( l_42 [6270] & !i[1820]) | ( l_42 [6271] &  i[1820]);
assign l_41[5185]    = ( l_42 [6272] & !i[1820]) | ( l_42 [6273] &  i[1820]);
assign l_41[5186]    = ( l_42 [6274] & !i[1820]) | ( l_42 [6275] &  i[1820]);
assign l_41[5187]    = ( l_42 [6276] & !i[1820]) | ( l_42 [6277] &  i[1820]);
assign l_41[5188]    = ( l_42 [6278] & !i[1820]) | ( l_42 [6279] &  i[1820]);
assign l_41[5189]    = ( l_42 [6280] & !i[1820]) | ( l_42 [6281] &  i[1820]);
assign l_41[5190]    = ( l_42 [6282] & !i[1820]) | ( l_42 [6283] &  i[1820]);
assign l_41[5191]    = ( l_42 [6284] & !i[1820]) | ( l_42 [6285] &  i[1820]);
assign l_41[5192]    = ( l_42 [6286] & !i[1820]) | ( l_42 [6287] &  i[1820]);
assign l_41[5193]    = ( l_42 [6288] & !i[1820]) | ( l_42 [6289] &  i[1820]);
assign l_41[5194]    = ( l_42 [6290] & !i[1820]) | ( l_42 [6291] &  i[1820]);
assign l_41[5195]    = ( l_42 [6292] & !i[1820]) | ( l_42 [6293] &  i[1820]);
assign l_41[5196]    = ( l_42 [6294] & !i[1820]) | ( l_42 [6295] &  i[1820]);
assign l_41[5197]    = ( l_42 [6296] & !i[1820]) | ( l_42 [6297] &  i[1820]);
assign l_41[5198]    = ( l_42 [6298] & !i[1820]) | ( l_42 [6299] &  i[1820]);
assign l_41[5199]    = ( l_42 [6300] & !i[1820]) | ( l_42 [6301] &  i[1820]);
assign l_41[5200]    = ( l_42 [6302] & !i[1820]) | ( l_42 [6303] &  i[1820]);
assign l_41[5201]    = ( l_42 [6304] & !i[1820]) | ( l_42 [6305] &  i[1820]);
assign l_41[5202]    = ( l_42 [6306] & !i[1820]) | ( l_42 [6307] &  i[1820]);
assign l_41[5203]    = ( l_42 [6308] & !i[1820]) | ( l_42 [6309] &  i[1820]);
assign l_41[5204]    = ( l_42 [6310] & !i[1820]) | ( l_42 [6311] &  i[1820]);
assign l_41[5205]    = ( l_42 [6312] & !i[1820]) | ( l_42 [6313] &  i[1820]);
assign l_41[5206]    = ( l_42 [6314] & !i[1820]) | ( l_42 [6315] &  i[1820]);
assign l_41[5207]    = ( l_42 [6316] & !i[1820]) | ( l_42 [6317] &  i[1820]);
assign l_41[5208]    = ( l_42 [6318] & !i[1820]) | ( l_42 [6319] &  i[1820]);
assign l_41[5209]    = ( l_42 [6320] & !i[1820]) | ( l_42 [6321] &  i[1820]);
assign l_41[5210]    = ( l_42 [6322] & !i[1820]) | ( l_42 [6323] &  i[1820]);
assign l_41[5211]    = ( l_42 [6324] & !i[1820]) | ( l_42 [6325] &  i[1820]);
assign l_41[5212]    = ( l_42 [6326] & !i[1820]) | ( l_42 [6327] &  i[1820]);
assign l_41[5213]    = ( l_42 [6328] & !i[1820]) | ( l_42 [6329] &  i[1820]);
assign l_41[5214]    = ( l_42 [6330] & !i[1820]) | ( l_42 [6331] &  i[1820]);
assign l_41[5215]    = ( l_42 [6332] & !i[1820]) | ( l_42 [6333] &  i[1820]);
assign l_41[5216]    = ( l_42 [6334] & !i[1820]) | ( l_42 [6335] &  i[1820]);
assign l_41[5217]    = ( l_42 [6336] & !i[1820]) | ( l_42 [6337] &  i[1820]);
assign l_41[5218]    = ( l_42 [6338] & !i[1820]) | ( l_42 [6339] &  i[1820]);
assign l_41[5219]    = ( l_42 [6340] & !i[1820]) | ( l_42 [6341] &  i[1820]);
assign l_41[5220]    = ( l_42 [6342] & !i[1820]) | ( l_42 [6343] &  i[1820]);
assign l_41[5221]    = ( l_42 [6344] & !i[1820]) | ( l_42 [6345] &  i[1820]);
assign l_41[5222]    = ( l_42 [6346] & !i[1820]) | ( l_42 [6347] &  i[1820]);
assign l_41[5223]    = ( l_42 [6348] & !i[1820]) | ( l_42 [6349] &  i[1820]);
assign l_41[5224]    = ( l_42 [6350] & !i[1820]) | ( l_42 [6351] &  i[1820]);
assign l_41[5225]    = ( l_42 [6352] & !i[1820]) | ( l_42 [6353] &  i[1820]);
assign l_41[5226]    = ( l_42 [6354] & !i[1820]) | ( l_42 [6355] &  i[1820]);
assign l_41[5227]    = ( l_42 [6356] & !i[1820]) | ( l_42 [6357] &  i[1820]);
assign l_41[5228]    = ( l_42 [6358] & !i[1820]) | ( l_42 [6359] &  i[1820]);
assign l_41[5229]    = ( l_42 [6360] & !i[1820]) | ( l_42 [6361] &  i[1820]);
assign l_41[5230]    = ( l_42 [6362] & !i[1820]) | ( l_42 [6363] &  i[1820]);
assign l_41[5231]    = ( l_42 [6364] & !i[1820]) | ( l_42 [6365] &  i[1820]);
assign l_41[5232]    = ( l_42 [6366] & !i[1820]) | ( l_42 [6367] &  i[1820]);
assign l_41[5233]    = ( l_42 [6368] & !i[1820]) | ( l_42 [6369] &  i[1820]);
assign l_41[5234]    = ( l_42 [6370] & !i[1820]) | ( l_42 [6371] &  i[1820]);
assign l_41[5235]    = ( l_42 [6372] & !i[1820]) | ( l_42 [6373] &  i[1820]);
assign l_41[5236]    = ( l_42 [6374] & !i[1820]) | ( l_42 [6375] &  i[1820]);
assign l_41[5237]    = ( l_42 [6376] & !i[1820]) | ( l_42 [6377] &  i[1820]);
assign l_41[5238]    = ( l_42 [6378] & !i[1820]) | ( l_42 [6379] &  i[1820]);
assign l_41[5239]    = ( l_42 [6380] & !i[1820]) | ( l_42 [6381] &  i[1820]);
assign l_41[5240]    = ( l_42 [6382] & !i[1820]) | ( l_42 [6383] &  i[1820]);
assign l_41[5241]    = ( l_42 [6384] & !i[1820]) | ( l_42 [6385] &  i[1820]);
assign l_41[5242]    = ( l_42 [6386] & !i[1820]) | ( l_42 [6387] &  i[1820]);
assign l_41[5243]    = ( l_42 [6388] & !i[1820]) | ( l_42 [6389] &  i[1820]);
assign l_41[5244]    = ( l_42 [6390] & !i[1820]) | ( l_42 [6391] &  i[1820]);
assign l_41[5245]    = ( l_42 [6392] & !i[1820]) | ( l_42 [6393] &  i[1820]);
assign l_41[5246]    = ( l_42 [6394] & !i[1820]) | ( l_42 [6395] &  i[1820]);
assign l_41[5247]    = ( l_42 [6396] & !i[1820]) | ( l_42 [6397] &  i[1820]);
assign l_41[5248]    = ( l_42 [6398] & !i[1820]) | ( l_42 [6399] &  i[1820]);
assign l_41[5249]    = ( l_42 [6400] & !i[1820]) | ( l_42 [6401] &  i[1820]);
assign l_41[5250]    = ( l_42 [6402] & !i[1820]) | ( l_42 [6403] &  i[1820]);
assign l_41[5251]    = ( l_42 [6404] & !i[1820]) | ( l_42 [6405] &  i[1820]);
assign l_41[5252]    = ( l_42 [6406] & !i[1820]) | ( l_42 [6407] &  i[1820]);
assign l_41[5253]    = ( l_42 [6408] & !i[1820]) | ( l_42 [6409] &  i[1820]);
assign l_41[5254]    = ( l_42 [6410] & !i[1820]) | ( l_42 [6411] &  i[1820]);
assign l_41[5255]    = ( l_42 [6412] & !i[1820]) | ( l_42 [6413] &  i[1820]);
assign l_41[5256]    = ( l_42 [6414] & !i[1820]) | ( l_42 [6415] &  i[1820]);
assign l_41[5257]    = ( l_42 [6416] & !i[1820]) | ( l_42 [6417] &  i[1820]);
assign l_41[5258]    = ( l_42 [6418] & !i[1820]) | ( l_42 [6419] &  i[1820]);
assign l_41[5259]    = ( l_42 [6420] & !i[1820]) | ( l_42 [6421] &  i[1820]);
assign l_41[5260]    = ( l_42 [6422] & !i[1820]) | ( l_42 [6423] &  i[1820]);
assign l_41[5261]    = ( l_42 [6424] & !i[1820]) | ( l_42 [6425] &  i[1820]);
assign l_41[5262]    = ( l_42 [6426] & !i[1820]) | ( l_42 [6427] &  i[1820]);
assign l_41[5263]    = ( l_42 [6428] & !i[1820]) | ( l_42 [6429] &  i[1820]);
assign l_41[5264]    = ( l_42 [6430] & !i[1820]) | ( l_42 [6431] &  i[1820]);
assign l_41[5265]    = ( l_42 [6432] & !i[1820]) | ( l_42 [6433] &  i[1820]);
assign l_41[5266]    = ( l_42 [6434] & !i[1820]) | ( l_42 [6435] &  i[1820]);
assign l_41[5267]    = ( l_42 [6436] & !i[1820]) | ( l_42 [6437] &  i[1820]);
assign l_41[5268]    = ( l_42 [6438] & !i[1820]) | ( l_42 [6439] &  i[1820]);
assign l_41[5269]    = ( l_42 [6440] & !i[1820]) | ( l_42 [6441] &  i[1820]);
assign l_41[5270]    = ( l_42 [6442] & !i[1820]) | ( l_42 [6443] &  i[1820]);
assign l_41[5271]    = ( l_42 [6444] & !i[1820]) | ( l_42 [6445] &  i[1820]);
assign l_41[5272]    = ( l_42 [6446] & !i[1820]) | ( l_42 [6447] &  i[1820]);
assign l_41[5273]    = ( l_42 [6448] & !i[1820]) | ( l_42 [6449] &  i[1820]);
assign l_41[5274]    = ( l_42 [6450] & !i[1820]) | ( l_42 [6451] &  i[1820]);
assign l_41[5275]    = ( l_42 [6452] & !i[1820]) | ( l_42 [6453] &  i[1820]);
assign l_41[5276]    = ( l_42 [6454] & !i[1820]) | ( l_42 [6455] &  i[1820]);
assign l_41[5277]    = ( l_42 [6456] & !i[1820]) | ( l_42 [6457] &  i[1820]);
assign l_41[5278]    = ( l_42 [6458] & !i[1820]) | ( l_42 [6459] &  i[1820]);
assign l_41[5279]    = ( l_42 [6460] & !i[1820]) | ( l_42 [6461] &  i[1820]);
assign l_41[5280]    = ( l_42 [6462] & !i[1820]) | ( l_42 [6463] &  i[1820]);
assign l_41[5281]    = ( l_42 [6464] & !i[1820]) | ( l_42 [6465] &  i[1820]);
assign l_41[5282]    = ( l_42 [6466] & !i[1820]) | ( l_42 [6467] &  i[1820]);
assign l_41[5283]    = ( l_42 [6468] & !i[1820]) | ( l_42 [6469] &  i[1820]);
assign l_41[5284]    = ( l_42 [6470] & !i[1820]) | ( l_42 [6471] &  i[1820]);
assign l_41[5285]    = ( l_42 [6472] & !i[1820]) | ( l_42 [6473] &  i[1820]);
assign l_41[5286]    = ( l_42 [6474] & !i[1820]) | ( l_42 [6475] &  i[1820]);
assign l_41[5287]    = ( l_42 [6476] & !i[1820]) | ( l_42 [6477] &  i[1820]);
assign l_41[5288]    = ( l_42 [6478] & !i[1820]) | ( l_42 [6479] &  i[1820]);
assign l_41[5289]    = ( l_42 [6480] & !i[1820]) | ( l_42 [6481] &  i[1820]);
assign l_41[5290]    = ( l_42 [6482] & !i[1820]) | ( l_42 [6483] &  i[1820]);
assign l_41[5291]    = ( l_42 [6484] & !i[1820]) | ( l_42 [6485] &  i[1820]);
assign l_41[5292]    = ( l_42 [6486] & !i[1820]) | ( l_42 [6487] &  i[1820]);
assign l_41[5293]    = ( l_42 [6488] & !i[1820]) | ( l_42 [6489] &  i[1820]);
assign l_41[5294]    = ( l_42 [6490] & !i[1820]) | ( l_42 [6491] &  i[1820]);
assign l_41[5295]    = ( l_42 [6492] & !i[1820]) | ( l_42 [6493] &  i[1820]);
assign l_41[5296]    = ( l_42 [6494] & !i[1820]) | ( l_42 [6495] &  i[1820]);
assign l_41[5297]    = ( l_42 [6496] & !i[1820]) | ( l_42 [6497] &  i[1820]);
assign l_41[5298]    = ( l_42 [6498] & !i[1820]) | ( l_42 [6499] &  i[1820]);
assign l_41[5299]    = ( l_42 [6500] & !i[1820]) | ( l_42 [6501] &  i[1820]);
assign l_41[5300]    = ( l_42 [6502] & !i[1820]) | ( l_42 [6503] &  i[1820]);
assign l_41[5301]    = ( l_42 [6504] & !i[1820]) | ( l_42 [6505] &  i[1820]);
assign l_41[5302]    = ( l_42 [6506] & !i[1820]) | ( l_42 [6507] &  i[1820]);
assign l_41[5303]    = ( l_42 [6508] & !i[1820]) | ( l_42 [6509] &  i[1820]);
assign l_41[5304]    = ( l_42 [6510] & !i[1820]) | ( l_42 [6511] &  i[1820]);
assign l_41[5305]    = ( l_42 [6512] & !i[1820]) | ( l_42 [6513] &  i[1820]);
assign l_41[5306]    = ( l_42 [6514] & !i[1820]) | ( l_42 [6515] &  i[1820]);
assign l_41[5307]    = ( l_42 [6516] & !i[1820]) | ( l_42 [6517] &  i[1820]);
assign l_41[5308]    = ( l_42 [6518] & !i[1820]) | ( l_42 [6519] &  i[1820]);
assign l_41[5309]    = ( l_42 [6520] & !i[1820]) | ( l_42 [6521] &  i[1820]);
assign l_41[5310]    = ( l_42 [6522] & !i[1820]) | ( l_42 [6523] &  i[1820]);
assign l_41[5311]    = ( l_42 [6524] & !i[1820]) | ( l_42 [6525] &  i[1820]);
assign l_41[5312]    = ( l_42 [6526] & !i[1820]) | ( l_42 [6527] &  i[1820]);
assign l_41[5313]    = ( l_42 [6528] & !i[1820]) | ( l_42 [6529] &  i[1820]);
assign l_41[5314]    = ( l_42 [6530] & !i[1820]) | ( l_42 [6531] &  i[1820]);
assign l_41[5315]    = ( l_42 [6532] & !i[1820]) | ( l_42 [6533] &  i[1820]);
assign l_41[5316]    = ( l_42 [6534] & !i[1820]) | ( l_42 [6535] &  i[1820]);
assign l_41[5317]    = ( l_42 [6536] & !i[1820]) | ( l_42 [6537] &  i[1820]);
assign l_41[5318]    = ( l_42 [6538] & !i[1820]) | ( l_42 [6539] &  i[1820]);
assign l_41[5319]    = ( l_42 [6540] & !i[1820]) | ( l_42 [6541] &  i[1820]);
assign l_41[5320]    = ( l_42 [6542] & !i[1820]) | ( l_42 [6543] &  i[1820]);
assign l_41[5321]    = ( l_42 [6544] & !i[1820]) | ( l_42 [6545] &  i[1820]);
assign l_41[5322]    = ( l_42 [6546] & !i[1820]) | ( l_42 [6547] &  i[1820]);
assign l_41[5323]    = ( l_42 [6548] & !i[1820]) | ( l_42 [6549] &  i[1820]);
assign l_41[5324]    = ( l_42 [6550] & !i[1820]) | ( l_42 [6551] &  i[1820]);
assign l_41[5325]    = ( l_42 [6552] & !i[1820]) | ( l_42 [6553] &  i[1820]);
assign l_41[5326]    = ( l_42 [6554] & !i[1820]) | ( l_42 [6555] &  i[1820]);
assign l_41[5327]    = ( l_42 [6556] & !i[1820]) | ( l_42 [6557] &  i[1820]);
assign l_41[5328]    = ( l_42 [6558] & !i[1820]) | ( l_42 [6559] &  i[1820]);
assign l_41[5329]    = ( l_42 [6560] & !i[1820]) | ( l_42 [6561] &  i[1820]);
assign l_41[5330]    = ( l_42 [6562] & !i[1820]) | ( l_42 [6563] &  i[1820]);
assign l_41[5331]    = ( l_42 [6564] & !i[1820]) | ( l_42 [6565] &  i[1820]);
assign l_41[5332]    = ( l_42 [6566] & !i[1820]) | ( l_42 [6567] &  i[1820]);
assign l_41[5333]    = ( l_42 [6568] & !i[1820]) | ( l_42 [6569] &  i[1820]);
assign l_41[5334]    = ( l_42 [6570] & !i[1820]) | ( l_42 [6571] &  i[1820]);
assign l_41[5335]    = ( l_42 [6572] & !i[1820]) | ( l_42 [6573] &  i[1820]);
assign l_41[5336]    = ( l_42 [6574] & !i[1820]) | ( l_42 [6575] &  i[1820]);
assign l_41[5337]    = ( l_42 [6576] & !i[1820]) | ( l_42 [6577] &  i[1820]);
assign l_41[5338]    = ( l_42 [6578] & !i[1820]) | ( l_42 [6579] &  i[1820]);
assign l_41[5339]    = ( l_42 [6580] & !i[1820]) | ( l_42 [6581] &  i[1820]);
assign l_41[5340]    = ( l_42 [6582] & !i[1820]) | ( l_42 [6583] &  i[1820]);
assign l_41[5341]    = ( l_42 [6584] & !i[1820]) | ( l_42 [6585] &  i[1820]);
assign l_41[5342]    = ( l_42 [6586] & !i[1820]) | ( l_42 [6587] &  i[1820]);
assign l_41[5343]    = ( l_42 [6588] & !i[1820]) | ( l_42 [6589] &  i[1820]);
assign l_41[5344]    = ( l_42 [6590] & !i[1820]) | ( l_42 [6591] &  i[1820]);
assign l_41[5345]    = ( l_42 [6592] & !i[1820]) | ( l_42 [6593] &  i[1820]);
assign l_41[5346]    = ( l_42 [6594] & !i[1820]) | ( l_42 [6595] &  i[1820]);
assign l_41[5347]    = ( l_42 [6596] & !i[1820]) | ( l_42 [6597] &  i[1820]);
assign l_41[5348]    = ( l_42 [6598] & !i[1820]) | ( l_42 [6599] &  i[1820]);
assign l_41[5349]    = ( l_42 [6600] & !i[1820]) | ( l_42 [6601] &  i[1820]);
assign l_41[5350]    = ( l_42 [6602] & !i[1820]) | ( l_42 [6603] &  i[1820]);
assign l_41[5351]    = ( l_42 [6604] & !i[1820]) | ( l_42 [6605] &  i[1820]);
assign l_41[5352]    = ( l_42 [6606] & !i[1820]) | ( l_42 [6607] &  i[1820]);
assign l_41[5353]    = ( l_42 [6608] & !i[1820]) | ( l_42 [6609] &  i[1820]);
assign l_41[5354]    = ( l_42 [6610] & !i[1820]) | ( l_42 [6611] &  i[1820]);
assign l_41[5355]    = ( l_42 [6612] & !i[1820]) | ( l_42 [6613] &  i[1820]);
assign l_41[5356]    = ( l_42 [6614] & !i[1820]) | ( l_42 [6615] &  i[1820]);
assign l_41[5357]    = ( l_42 [6616] & !i[1820]) | ( l_42 [6617] &  i[1820]);
assign l_41[5358]    = ( l_42 [6618] & !i[1820]) | ( l_42 [6619] &  i[1820]);
assign l_41[5359]    = ( l_42 [6620] & !i[1820]) | ( l_42 [6621] &  i[1820]);
assign l_41[5360]    = ( l_42 [6622] & !i[1820]) | ( l_42 [6623] &  i[1820]);
assign l_41[5361]    = ( l_42 [6624] & !i[1820]) | ( l_42 [6625] &  i[1820]);
assign l_41[5362]    = ( l_42 [6626] & !i[1820]) | ( l_42 [6627] &  i[1820]);
assign l_41[5363]    = ( l_42 [6628] & !i[1820]) | ( l_42 [6629] &  i[1820]);
assign l_41[5364]    = ( l_42 [6630] & !i[1820]) | ( l_42 [6631] &  i[1820]);
assign l_41[5365]    = ( l_42 [6632] & !i[1820]) | ( l_42 [6633] &  i[1820]);
assign l_41[5366]    = ( l_42 [6634] & !i[1820]) | ( l_42 [6635] &  i[1820]);
assign l_41[5367]    = ( l_42 [6636] & !i[1820]) | ( l_42 [6637] &  i[1820]);
assign l_41[5368]    = ( l_42 [6638] & !i[1820]) | ( l_42 [6639] &  i[1820]);
assign l_41[5369]    = ( l_42 [6640] & !i[1820]) | ( l_42 [6641] &  i[1820]);
assign l_41[5370]    = ( l_42 [6642] & !i[1820]) | ( l_42 [6643] &  i[1820]);
assign l_41[5371]    = ( l_42 [6644] & !i[1820]) | ( l_42 [6645] &  i[1820]);
assign l_41[5372]    = ( l_42 [6646] & !i[1820]) | ( l_42 [6647] &  i[1820]);
assign l_41[5373]    = ( l_42 [6648] & !i[1820]) | ( l_42 [6649] &  i[1820]);
assign l_41[5374]    = ( l_42 [6650] & !i[1820]) | ( l_42 [6651] &  i[1820]);
assign l_41[5375]    = ( l_42 [6652] & !i[1820]) | ( l_42 [6653] &  i[1820]);
assign l_41[5376]    = ( l_42 [6654] & !i[1820]) | ( l_42 [6655] &  i[1820]);
assign l_41[5377]    = ( l_42 [6656] & !i[1820]) | ( l_42 [6657] &  i[1820]);
assign l_41[5378]    = ( l_42 [6658] & !i[1820]) | ( l_42 [6659] &  i[1820]);
assign l_41[5379]    = ( l_42 [6660] & !i[1820]) | ( l_42 [6661] &  i[1820]);
assign l_41[5380]    = ( l_42 [6662] & !i[1820]) | ( l_42 [6663] &  i[1820]);
assign l_41[5381]    = ( l_42 [6664] & !i[1820]) | ( l_42 [6665] &  i[1820]);
assign l_41[5382]    = ( l_42 [6666] & !i[1820]) | ( l_42 [6667] &  i[1820]);
assign l_41[5383]    = ( l_42 [6668] & !i[1820]) | ( l_42 [6669] &  i[1820]);
assign l_41[5384]    = ( l_42 [6670] & !i[1820]) | ( l_42 [6671] &  i[1820]);
assign l_41[5385]    = ( l_42 [6672] & !i[1820]) | ( l_42 [6673] &  i[1820]);
assign l_41[5386]    = ( l_42 [6674] & !i[1820]) | ( l_42 [6675] &  i[1820]);
assign l_41[5387]    = ( l_42 [6676] & !i[1820]) | ( l_42 [6677] &  i[1820]);
assign l_41[5388]    = ( l_42 [6678] & !i[1820]) | ( l_42 [6679] &  i[1820]);
assign l_41[5389]    = ( l_42 [6680] & !i[1820]) | ( l_42 [6681] &  i[1820]);
assign l_41[5390]    = ( l_42 [6682] & !i[1820]) | ( l_42 [6683] &  i[1820]);
assign l_41[5391]    = ( l_42 [6684] & !i[1820]) | ( l_42 [6685] &  i[1820]);
assign l_41[5392]    = ( l_42 [6686] & !i[1820]) | ( l_42 [6687] &  i[1820]);
assign l_41[5393]    = ( l_42 [6688] & !i[1820]) | ( l_42 [6689] &  i[1820]);
assign l_41[5394]    = ( l_42 [6690] & !i[1820]) | ( l_42 [6691] &  i[1820]);
assign l_41[5395]    = ( l_42 [6692] & !i[1820]) | ( l_42 [6693] &  i[1820]);
assign l_41[5396]    = ( l_42 [6694] & !i[1820]) | ( l_42 [6695] &  i[1820]);
assign l_41[5397]    = ( l_42 [6696] & !i[1820]) | ( l_42 [6697] &  i[1820]);
assign l_41[5398]    = ( l_42 [6698] & !i[1820]) | ( l_42 [6699] &  i[1820]);
assign l_41[5399]    = ( l_42 [6700] & !i[1820]) | ( l_42 [6701] &  i[1820]);
assign l_41[5400]    = ( l_42 [6702] & !i[1820]) | ( l_42 [6703] &  i[1820]);
assign l_41[5401]    = ( l_42 [6704] & !i[1820]) | ( l_42 [6705] &  i[1820]);
assign l_41[5402]    = ( l_42 [6706] & !i[1820]) | ( l_42 [6707] &  i[1820]);
assign l_41[5403]    = ( l_42 [6708] & !i[1820]) | ( l_42 [6709] &  i[1820]);
assign l_41[5404]    = ( l_42 [6710] & !i[1820]) | ( l_42 [6711] &  i[1820]);
assign l_41[5405]    = ( l_42 [6712] & !i[1820]) | ( l_42 [6713] &  i[1820]);
assign l_41[5406]    = ( l_42 [6714] & !i[1820]) | ( l_42 [6715] &  i[1820]);
assign l_41[5407]    = ( l_42 [6716] & !i[1820]) | ( l_42 [6717] &  i[1820]);
assign l_41[5408]    = ( l_42 [6718] & !i[1820]) | ( l_42 [6719] &  i[1820]);
assign l_41[5409]    = ( l_42 [6720] & !i[1820]) | ( l_42 [6721] &  i[1820]);
assign l_41[5410]    = ( l_42 [6722] & !i[1820]) | ( l_42 [6723] &  i[1820]);
assign l_41[5411]    = ( l_42 [6724] & !i[1820]) | ( l_42 [6725] &  i[1820]);
assign l_41[5412]    = ( l_42 [6726] & !i[1820]) | ( l_42 [6727] &  i[1820]);
assign l_41[5413]    = ( l_42 [6728] & !i[1820]) | ( l_42 [6729] &  i[1820]);
assign l_41[5414]    = ( l_42 [6730] & !i[1820]) | ( l_42 [6731] &  i[1820]);
assign l_41[5415]    = ( l_42 [6732] & !i[1820]) | ( l_42 [6733] &  i[1820]);
assign l_41[5416]    = ( l_42 [6734] & !i[1820]) | ( l_42 [6735] &  i[1820]);
assign l_41[5417]    = ( l_42 [6736] & !i[1820]) | ( l_42 [6737] &  i[1820]);
assign l_41[5418]    = ( l_42 [6738] & !i[1820]) | ( l_42 [6739] &  i[1820]);
assign l_41[5419]    = ( l_42 [6740] & !i[1820]) | ( l_42 [6741] &  i[1820]);
assign l_41[5420]    = ( l_42 [6742] & !i[1820]) | ( l_42 [6743] &  i[1820]);
assign l_41[5421]    = ( l_42 [6744] & !i[1820]) | ( l_42 [6745] &  i[1820]);
assign l_41[5422]    = ( l_42 [6746] & !i[1820]) | ( l_42 [6747] &  i[1820]);
assign l_41[5423]    = ( l_42 [6748] & !i[1820]) | ( l_42 [6749] &  i[1820]);
assign l_41[5424]    = ( l_42 [6750] & !i[1820]) | ( l_42 [6751] &  i[1820]);
assign l_41[5425]    = ( l_42 [6752] & !i[1820]) | ( l_42 [6753] &  i[1820]);
assign l_41[5426]    = ( l_42 [6754] & !i[1820]) | ( l_42 [6755] &  i[1820]);
assign l_41[5427]    = ( l_42 [6756] & !i[1820]) | ( l_42 [6757] &  i[1820]);
assign l_41[5428]    = ( l_42 [6758] & !i[1820]) | ( l_42 [6759] &  i[1820]);
assign l_41[5429]    = ( l_42 [6760] & !i[1820]) | ( l_42 [6761] &  i[1820]);
assign l_41[5430]    = ( l_42 [6762] & !i[1820]) | ( l_42 [6763] &  i[1820]);
assign l_41[5431]    = ( l_42 [6764] & !i[1820]) | ( l_42 [6765] &  i[1820]);
assign l_41[5432]    = ( l_42 [6766] & !i[1820]) | ( l_42 [6767] &  i[1820]);
assign l_41[5433]    = ( l_42 [6768] & !i[1820]) | ( l_42 [6769] &  i[1820]);
assign l_41[5434]    = ( l_42 [6770] & !i[1820]) | ( l_42 [6771] &  i[1820]);
assign l_41[5435]    = ( l_42 [6772] & !i[1820]) | ( l_42 [6773] &  i[1820]);
assign l_41[5436]    = ( l_42 [6774] & !i[1820]) | ( l_42 [6775] &  i[1820]);
assign l_41[5437]    = ( l_42 [6776] & !i[1820]) | ( l_42 [6777] &  i[1820]);
assign l_41[5438]    = ( l_42 [6778] & !i[1820]) | ( l_42 [6779] &  i[1820]);
assign l_41[5439]    = ( l_42 [6780] & !i[1820]) | ( l_42 [6781] &  i[1820]);
assign l_41[5440]    = ( l_42 [6782] & !i[1820]) | ( l_42 [6783] &  i[1820]);
assign l_41[5441]    = ( l_42 [6784] & !i[1820]) | ( l_42 [6785] &  i[1820]);
assign l_41[5442]    = ( l_42 [6786] & !i[1820]) | ( l_42 [6787] &  i[1820]);
assign l_41[5443]    = ( l_42 [6788] & !i[1820]) | ( l_42 [6789] &  i[1820]);
assign l_41[5444]    = ( l_42 [6790] & !i[1820]) | ( l_42 [6791] &  i[1820]);
assign l_41[5445]    = ( l_42 [6792] & !i[1820]) | ( l_42 [6793] &  i[1820]);
assign l_41[5446]    = ( l_42 [6794] & !i[1820]) | ( l_42 [6795] &  i[1820]);
assign l_41[5447]    = ( l_42 [6796] & !i[1820]) | ( l_42 [6797] &  i[1820]);
assign l_41[5448]    = ( l_42 [6798] & !i[1820]) | ( l_42 [6799] &  i[1820]);
assign l_41[5449]    = ( l_42 [6800] & !i[1820]) | ( l_42 [6801] &  i[1820]);
assign l_41[5450]    = ( l_42 [6802] & !i[1820]) | ( l_42 [6803] &  i[1820]);
assign l_41[5451]    = ( l_42 [6804] & !i[1820]) | ( l_42 [6805] &  i[1820]);
assign l_41[5452]    = ( l_42 [6806] & !i[1820]) | ( l_42 [6807] &  i[1820]);
assign l_41[5453]    = ( l_42 [6808] & !i[1820]) | ( l_42 [6809] &  i[1820]);
assign l_41[5454]    = ( l_42 [6810] & !i[1820]) | ( l_42 [6811] &  i[1820]);
assign l_41[5455]    = ( l_42 [6812] & !i[1820]) | ( l_42 [6813] &  i[1820]);
assign l_41[5456]    = ( l_42 [6814] & !i[1820]) | ( l_42 [6815] &  i[1820]);
assign l_41[5457]    = ( l_42 [6816] & !i[1820]) | ( l_42 [6817] &  i[1820]);
assign l_41[5458]    = ( l_42 [6818] & !i[1820]) | ( l_42 [6819] &  i[1820]);
assign l_41[5459]    = ( l_42 [6820] & !i[1820]) | ( l_42 [6821] &  i[1820]);
assign l_41[5460]    = ( l_42 [6822] & !i[1820]) | ( l_42 [6823] &  i[1820]);
assign l_41[5461]    = ( l_42 [6824] & !i[1820]) | ( l_42 [6825] &  i[1820]);
assign l_41[5462]    = ( l_42 [6826] & !i[1820]) | ( l_42 [6827] &  i[1820]);
assign l_41[5463]    = ( l_42 [6828] & !i[1820]) | ( l_42 [6829] &  i[1820]);
assign l_41[5464]    = ( l_42 [6830] & !i[1820]) | ( l_42 [6831] &  i[1820]);
assign l_41[5465]    = ( l_42 [6832] & !i[1820]) | ( l_42 [6833] &  i[1820]);
assign l_41[5466]    = ( l_42 [6834] & !i[1820]) | ( l_42 [6835] &  i[1820]);
assign l_41[5467]    = ( l_42 [6836] & !i[1820]) | ( l_42 [6837] &  i[1820]);
assign l_41[5468]    = ( l_42 [6838] & !i[1820]) | ( l_42 [6839] &  i[1820]);
assign l_41[5469]    = ( l_42 [6840] & !i[1820]) | ( l_42 [6841] &  i[1820]);
assign l_41[5470]    = ( l_42 [6842] & !i[1820]) | ( l_42 [6843] &  i[1820]);
assign l_41[5471]    = ( l_42 [6844] & !i[1820]) | ( l_42 [6845] &  i[1820]);
assign l_41[5472]    = ( l_42 [6846] & !i[1820]) | ( l_42 [6847] &  i[1820]);
assign l_41[5473]    = ( l_42 [6848] & !i[1820]) | ( l_42 [6849] &  i[1820]);
assign l_41[5474]    = ( l_42 [6850] & !i[1820]) | ( l_42 [6851] &  i[1820]);
assign l_41[5475]    = ( l_42 [6852] & !i[1820]) | ( l_42 [6853] &  i[1820]);
assign l_41[5476]    = ( l_42 [6854] & !i[1820]) | ( l_42 [6855] &  i[1820]);
assign l_41[5477]    = ( l_42 [6856] & !i[1820]) | ( l_42 [6857] &  i[1820]);
assign l_41[5478]    = ( l_42 [6858] & !i[1820]) | ( l_42 [6859] &  i[1820]);
assign l_41[5479]    = ( l_42 [6860] & !i[1820]) | ( l_42 [6861] &  i[1820]);
assign l_41[5480]    = ( l_42 [6862] & !i[1820]) | ( l_42 [6863] &  i[1820]);
assign l_41[5481]    = ( l_42 [6864] & !i[1820]) | ( l_42 [6865] &  i[1820]);
assign l_41[5482]    = ( l_42 [6866] & !i[1820]) | ( l_42 [6867] &  i[1820]);
assign l_41[5483]    = ( l_42 [6868] & !i[1820]) | ( l_42 [6869] &  i[1820]);
assign l_41[5484]    = ( l_42 [6870] & !i[1820]) | ( l_42 [6871] &  i[1820]);
assign l_41[5485]    = ( l_42 [6872] & !i[1820]) | ( l_42 [6873] &  i[1820]);
assign l_41[5486]    = ( l_42 [6874] & !i[1820]) | ( l_42 [6875] &  i[1820]);
assign l_41[5487]    = ( l_42 [6876] & !i[1820]) | ( l_42 [6877] &  i[1820]);
assign l_41[5488]    = ( l_42 [6878] & !i[1820]) | ( l_42 [6879] &  i[1820]);
assign l_41[5489]    = ( l_42 [6880] & !i[1820]) | ( l_42 [6881] &  i[1820]);
assign l_41[5490]    = ( l_42 [6882] & !i[1820]) | ( l_42 [6883] &  i[1820]);
assign l_41[5491]    = ( l_42 [6884] & !i[1820]) | ( l_42 [6885] &  i[1820]);
assign l_41[5492]    = ( l_42 [6886] & !i[1820]) | ( l_42 [6887] &  i[1820]);
assign l_41[5493]    = ( l_42 [6888] & !i[1820]) | ( l_42 [6889] &  i[1820]);
assign l_41[5494]    = ( l_42 [6890] & !i[1820]) | ( l_42 [6891] &  i[1820]);
assign l_41[5495]    = ( l_42 [6892] & !i[1820]) | ( l_42 [6893] &  i[1820]);
assign l_41[5496]    = ( l_42 [6894] & !i[1820]) | ( l_42 [6895] &  i[1820]);
assign l_41[5497]    = ( l_42 [6896] & !i[1820]) | ( l_42 [6897] &  i[1820]);
assign l_41[5498]    = ( l_42 [6898] & !i[1820]) | ( l_42 [6899] &  i[1820]);
assign l_41[5499]    = ( l_42 [6900] & !i[1820]) | ( l_42 [6901] &  i[1820]);
assign l_41[5500]    = ( l_42 [6902] & !i[1820]) | ( l_42 [6903] &  i[1820]);
assign l_41[5501]    = ( l_42 [6904] & !i[1820]) | ( l_42 [6905] &  i[1820]);
assign l_41[5502]    = ( l_42 [6906] & !i[1820]) | ( l_42 [6907] &  i[1820]);
assign l_41[5503]    = ( l_42 [6908] & !i[1820]) | ( l_42 [6909] &  i[1820]);
assign l_41[5504]    = ( l_42 [6910] & !i[1820]) | ( l_42 [6911] &  i[1820]);
assign l_41[5505]    = ( l_42 [6912] & !i[1820]) | ( l_42 [6913] &  i[1820]);
assign l_41[5506]    = ( l_42 [6914] & !i[1820]) | ( l_42 [6915] &  i[1820]);
assign l_41[5507]    = ( l_42 [6916] & !i[1820]) | ( l_42 [6917] &  i[1820]);
assign l_41[5508]    = ( l_42 [6918] & !i[1820]) | ( l_42 [6919] &  i[1820]);
assign l_41[5509]    = ( l_42 [6920] & !i[1820]) | ( l_42 [6921] &  i[1820]);
assign l_41[5510]    = ( l_42 [6922] & !i[1820]) | ( l_42 [6923] &  i[1820]);
assign l_41[5511]    = ( l_42 [6924] & !i[1820]) | ( l_42 [6925] &  i[1820]);
assign l_41[5512]    = ( l_42 [6926] & !i[1820]) | ( l_42 [6927] &  i[1820]);
assign l_41[5513]    = ( l_42 [6928] & !i[1820]) | ( l_42 [6929] &  i[1820]);
assign l_41[5514]    = ( l_42 [6930] & !i[1820]) | ( l_42 [6931] &  i[1820]);
assign l_41[5515]    = ( l_42 [6932] & !i[1820]) | ( l_42 [6933] &  i[1820]);
assign l_41[5516]    = ( l_42 [6934] & !i[1820]) | ( l_42 [6935] &  i[1820]);
assign l_41[5517]    = ( l_42 [6936] & !i[1820]) | ( l_42 [6937] &  i[1820]);
assign l_41[5518]    = ( l_42 [6938] & !i[1820]) | ( l_42 [6939] &  i[1820]);
assign l_41[5519]    = ( l_42 [6940] & !i[1820]) | ( l_42 [6941] &  i[1820]);
assign l_41[5520]    = ( l_42 [6942] & !i[1820]) | ( l_42 [6943] &  i[1820]);
assign l_41[5521]    = ( l_42 [6944] & !i[1820]) | ( l_42 [6945] &  i[1820]);
assign l_41[5522]    = ( l_42 [6946] & !i[1820]) | ( l_42 [6947] &  i[1820]);
assign l_41[5523]    = ( l_42 [6948] & !i[1820]) | ( l_42 [6949] &  i[1820]);
assign l_41[5524]    = ( l_42 [6950] & !i[1820]) | ( l_42 [6951] &  i[1820]);
assign l_41[5525]    = ( l_42 [6952] & !i[1820]) | ( l_42 [6953] &  i[1820]);
assign l_41[5526]    = ( l_42 [6954] & !i[1820]) | ( l_42 [6955] &  i[1820]);
assign l_41[5527]    = ( l_42 [6956] & !i[1820]) | ( l_42 [6957] &  i[1820]);
assign l_41[5528]    = ( l_42 [6958] & !i[1820]) | ( l_42 [6959] &  i[1820]);
assign l_41[5529]    = ( l_42 [6960] & !i[1820]) | ( l_42 [6961] &  i[1820]);
assign l_41[5530]    = ( l_42 [6962] & !i[1820]) | ( l_42 [6963] &  i[1820]);
assign l_41[5531]    = ( l_42 [6964] & !i[1820]) | ( l_42 [6965] &  i[1820]);
assign l_41[5532]    = ( l_42 [6966] & !i[1820]) | ( l_42 [6967] &  i[1820]);
assign l_41[5533]    = ( l_42 [6968] & !i[1820]) | ( l_42 [6969] &  i[1820]);
assign l_41[5534]    = ( l_42 [6970] & !i[1820]) | ( l_42 [6971] &  i[1820]);
assign l_41[5535]    = ( l_42 [6972] & !i[1820]) | ( l_42 [6973] &  i[1820]);
assign l_41[5536]    = ( l_42 [6974] & !i[1820]) | ( l_42 [6975] &  i[1820]);
assign l_41[5537]    = ( l_42 [6976] & !i[1820]) | ( l_42 [6977] &  i[1820]);
assign l_41[5538]    = ( l_42 [6978] & !i[1820]) | ( l_42 [6979] &  i[1820]);
assign l_41[5539]    = ( l_42 [6980] & !i[1820]) | ( l_42 [6981] &  i[1820]);
assign l_41[5540]    = ( l_42 [6982] & !i[1820]) | ( l_42 [6983] &  i[1820]);
assign l_41[5541]    = ( l_42 [6984] & !i[1820]) | ( l_42 [6985] &  i[1820]);
assign l_41[5542]    = ( l_42 [6986] & !i[1820]) | ( l_42 [6987] &  i[1820]);
assign l_41[5543]    = ( l_42 [6988] & !i[1820]) | ( l_42 [6989] &  i[1820]);
assign l_41[5544]    = ( l_42 [6990] & !i[1820]) | ( l_42 [6991] &  i[1820]);
assign l_41[5545]    = ( l_42 [6992] & !i[1820]) | ( l_42 [6993] &  i[1820]);
assign l_41[5546]    = ( l_42 [6994] & !i[1820]) | ( l_42 [6995] &  i[1820]);
assign l_41[5547]    = ( l_42 [6996] & !i[1820]) | ( l_42 [6997] &  i[1820]);
assign l_41[5548]    = ( l_42 [6998] & !i[1820]) | ( l_42 [6999] &  i[1820]);
assign l_41[5549]    = ( l_42 [7000] & !i[1820]) | ( l_42 [7001] &  i[1820]);
assign l_41[5550]    = ( l_42 [7002] & !i[1820]) | ( l_42 [7003] &  i[1820]);
assign l_41[5551]    = ( l_42 [7004] & !i[1820]) | ( l_42 [7005] &  i[1820]);
assign l_41[5552]    = ( l_42 [7006] & !i[1820]) | ( l_42 [7007] &  i[1820]);
assign l_41[5553]    = ( l_42 [7008] & !i[1820]) | ( l_42 [7009] &  i[1820]);
assign l_41[5554]    = ( l_42 [7010] & !i[1820]) | ( l_42 [7011] &  i[1820]);
assign l_41[5555]    = ( l_42 [7012] & !i[1820]) | ( l_42 [7013] &  i[1820]);
assign l_41[5556]    = ( l_42 [7014] & !i[1820]) | ( l_42 [7015] &  i[1820]);
assign l_41[5557]    = ( l_42 [7016] & !i[1820]) | ( l_42 [7017] &  i[1820]);
assign l_41[5558]    = ( l_42 [7018] & !i[1820]) | ( l_42 [7019] &  i[1820]);
assign l_41[5559]    = ( l_42 [7020] & !i[1820]) | ( l_42 [7021] &  i[1820]);
assign l_41[5560]    = ( l_42 [7022] & !i[1820]) | ( l_42 [7023] &  i[1820]);
assign l_41[5561]    = ( l_42 [7024] & !i[1820]) | ( l_42 [7025] &  i[1820]);
assign l_41[5562]    = ( l_42 [7026] & !i[1820]) | ( l_42 [7027] &  i[1820]);
assign l_41[5563]    = ( l_42 [7028] & !i[1820]) | ( l_42 [7029] &  i[1820]);
assign l_41[5564]    = ( l_42 [7030] & !i[1820]) | ( l_42 [7031] &  i[1820]);
assign l_41[5565]    = ( l_42 [7032] & !i[1820]) | ( l_42 [7033] &  i[1820]);
assign l_41[5566]    = ( l_42 [7034] & !i[1820]) | ( l_42 [7035] &  i[1820]);
assign l_41[5567]    = ( l_42 [7036] & !i[1820]) | ( l_42 [7037] &  i[1820]);
assign l_41[5568]    = ( l_42 [7038] & !i[1820]) | ( l_42 [7039] &  i[1820]);
assign l_41[5569]    = ( l_42 [7040] & !i[1820]) | ( l_42 [7041] &  i[1820]);
assign l_41[5570]    = ( l_42 [7042] & !i[1820]) | ( l_42 [7043] &  i[1820]);
assign l_41[5571]    = ( l_42 [7044] & !i[1820]) | ( l_42 [7045] &  i[1820]);
assign l_41[5572]    = ( l_42 [7046] & !i[1820]) | ( l_42 [7047] &  i[1820]);
assign l_41[5573]    = ( l_42 [7048] & !i[1820]) | ( l_42 [7049] &  i[1820]);
assign l_41[5574]    = ( l_42 [7050] & !i[1820]) | ( l_42 [7051] &  i[1820]);
assign l_41[5575]    = ( l_42 [7052] & !i[1820]) | ( l_42 [7053] &  i[1820]);
assign l_41[5576]    = ( l_42 [7054] & !i[1820]) | ( l_42 [7055] &  i[1820]);
assign l_41[5577]    = ( l_42 [7056] & !i[1820]) | ( l_42 [7057] &  i[1820]);
assign l_41[5578]    = ( l_42 [7058] & !i[1820]) | ( l_42 [7059] &  i[1820]);
assign l_41[5579]    = ( l_42 [7060] & !i[1820]) | ( l_42 [7061] &  i[1820]);
assign l_41[5580]    = ( l_42 [7062] & !i[1820]) | ( l_42 [7063] &  i[1820]);
assign l_41[5581]    = ( l_42 [7064] & !i[1820]) | ( l_42 [7065] &  i[1820]);
assign l_41[5582]    = ( l_42 [7066] & !i[1820]) | ( l_42 [7067] &  i[1820]);
assign l_41[5583]    = ( l_42 [7068] & !i[1820]) | ( l_42 [7069] &  i[1820]);
assign l_41[5584]    = ( l_42 [7070] & !i[1820]) | ( l_42 [7071] &  i[1820]);
assign l_41[5585]    = ( l_42 [7072] & !i[1820]) | ( l_42 [7073] &  i[1820]);
assign l_41[5586]    = ( l_42 [7074] & !i[1820]) | ( l_42 [7075] &  i[1820]);
assign l_41[5587]    = ( l_42 [7076] & !i[1820]) | ( l_42 [7077] &  i[1820]);
assign l_41[5588]    = ( l_42 [7078] & !i[1820]) | ( l_42 [7079] &  i[1820]);
assign l_41[5589]    = ( l_42 [7080] & !i[1820]) | ( l_42 [7081] &  i[1820]);
assign l_41[5590]    = ( l_42 [7082] & !i[1820]) | ( l_42 [7083] &  i[1820]);
assign l_41[5591]    = ( l_42 [7084] & !i[1820]) | ( l_42 [7085] &  i[1820]);
assign l_41[5592]    = ( l_42 [7086] & !i[1820]) | ( l_42 [7087] &  i[1820]);
assign l_41[5593]    = ( l_42 [7088] & !i[1820]) | ( l_42 [7089] &  i[1820]);
assign l_41[5594]    = ( l_42 [7090] & !i[1820]) | ( l_42 [7091] &  i[1820]);
assign l_41[5595]    = ( l_42 [7092] & !i[1820]) | ( l_42 [7093] &  i[1820]);
assign l_41[5596]    = ( l_42 [7094] & !i[1820]) | ( l_42 [7095] &  i[1820]);
assign l_41[5597]    = ( l_42 [7096] & !i[1820]) | ( l_42 [7097] &  i[1820]);
assign l_41[5598]    = ( l_42 [7098] & !i[1820]) | ( l_42 [7099] &  i[1820]);
assign l_41[5599]    = ( l_42 [7100] & !i[1820]) | ( l_42 [7101] &  i[1820]);
assign l_41[5600]    = ( l_42 [7102] & !i[1820]) | ( l_42 [7103] &  i[1820]);
assign l_41[5601]    = ( l_42 [7104] & !i[1820]) | ( l_42 [7105] &  i[1820]);
assign l_41[5602]    = ( l_42 [7106] & !i[1820]) | ( l_42 [7107] &  i[1820]);
assign l_41[5603]    = ( l_42 [7108] & !i[1820]) | ( l_42 [7109] &  i[1820]);
assign l_41[5604]    = ( l_42 [7110] & !i[1820]) | ( l_42 [7111] &  i[1820]);
assign l_41[5605]    = ( l_42 [7112] & !i[1820]) | ( l_42 [7113] &  i[1820]);
assign l_41[5606]    = ( l_42 [7114] & !i[1820]) | ( l_42 [7115] &  i[1820]);
assign l_41[5607]    = ( l_42 [7116] & !i[1820]) | ( l_42 [7117] &  i[1820]);
assign l_41[5608]    = ( l_42 [7118] & !i[1820]) | ( l_42 [7119] &  i[1820]);
assign l_41[5609]    = ( l_42 [7120] & !i[1820]) | ( l_42 [7121] &  i[1820]);
assign l_41[5610]    = ( l_42 [7122] & !i[1820]) | ( l_42 [7123] &  i[1820]);
assign l_41[5611]    = ( l_42 [7124] & !i[1820]) | ( l_42 [7125] &  i[1820]);
assign l_41[5612]    = ( l_42 [7126] & !i[1820]) | ( l_42 [7127] &  i[1820]);
assign l_41[5613]    = ( l_42 [7128] & !i[1820]) | ( l_42 [7129] &  i[1820]);
assign l_41[5614]    = ( l_42 [7130] & !i[1820]) | ( l_42 [7131] &  i[1820]);
assign l_41[5615]    = ( l_42 [7132] & !i[1820]) | ( l_42 [7133] &  i[1820]);
assign l_41[5616]    = ( l_42 [7134] & !i[1820]) | ( l_42 [7135] &  i[1820]);
assign l_41[5617]    = ( l_42 [7136] & !i[1820]) | ( l_42 [7137] &  i[1820]);
assign l_41[5618]    = ( l_42 [7138] & !i[1820]) | ( l_42 [7139] &  i[1820]);
assign l_41[5619]    = ( l_42 [7140] & !i[1820]) | ( l_42 [7141] &  i[1820]);
assign l_41[5620]    = ( l_42 [7142] & !i[1820]) | ( l_42 [7143] &  i[1820]);
assign l_41[5621]    = ( l_42 [7144] & !i[1820]) | ( l_42 [7145] &  i[1820]);
assign l_41[5622]    = ( l_42 [7146] & !i[1820]) | ( l_42 [7147] &  i[1820]);
assign l_41[5623]    = ( l_42 [7148] & !i[1820]) | ( l_42 [7149] &  i[1820]);
assign l_41[5624]    = ( l_42 [7150] & !i[1820]) | ( l_42 [7151] &  i[1820]);
assign l_41[5625]    = ( l_42 [7152] & !i[1820]) | ( l_42 [7153] &  i[1820]);
assign l_41[5626]    = ( l_42 [7154] & !i[1820]) | ( l_42 [7155] &  i[1820]);
assign l_41[5627]    = ( l_42 [7156] & !i[1820]) | ( l_42 [7157] &  i[1820]);
assign l_41[5628]    = ( l_42 [7158] & !i[1820]) | ( l_42 [7159] &  i[1820]);
assign l_41[5629]    = ( l_42 [7160] & !i[1820]) | ( l_42 [7161] &  i[1820]);
assign l_41[5630]    = ( l_42 [7162] & !i[1820]) | ( l_42 [7163] &  i[1820]);
assign l_41[5631]    = ( l_42 [7164] & !i[1820]) | ( l_42 [7165] &  i[1820]);
assign l_41[5632]    = ( l_42 [7166] & !i[1820]) | ( l_42 [7167] &  i[1820]);
assign l_41[5633]    = ( l_42 [7168] & !i[1820]) | ( l_42 [7169] &  i[1820]);
assign l_41[5634]    = ( l_42 [7170] & !i[1820]) | ( l_42 [7171] &  i[1820]);
assign l_41[5635]    = ( l_42 [7172] & !i[1820]) | ( l_42 [7173] &  i[1820]);
assign l_41[5636]    = ( l_42 [7174] & !i[1820]) | ( l_42 [7175] &  i[1820]);
assign l_41[5637]    = ( l_42 [7176] & !i[1820]) | ( l_42 [7177] &  i[1820]);
assign l_41[5638]    = ( l_42 [7178] & !i[1820]) | ( l_42 [7179] &  i[1820]);
assign l_41[5639]    = ( l_42 [7180] & !i[1820]) | ( l_42 [7181] &  i[1820]);
assign l_41[5640]    = ( l_42 [7182] & !i[1820]) | ( l_42 [7183] &  i[1820]);
assign l_41[5641]    = ( l_42 [7184] & !i[1820]) | ( l_42 [7185] &  i[1820]);
assign l_41[5642]    = ( l_42 [7186] & !i[1820]) | ( l_42 [7187] &  i[1820]);
assign l_41[5643]    = ( l_42 [7188] & !i[1820]) | ( l_42 [7189] &  i[1820]);
assign l_41[5644]    = ( l_42 [7190] & !i[1820]) | ( l_42 [7191] &  i[1820]);
assign l_41[5645]    = ( l_42 [7192] & !i[1820]) | ( l_42 [7193] &  i[1820]);
assign l_41[5646]    = ( l_42 [7194] & !i[1820]) | ( l_42 [7195] &  i[1820]);
assign l_41[5647]    = ( l_42 [7196] & !i[1820]) | ( l_42 [7197] &  i[1820]);
assign l_41[5648]    = ( l_42 [7198] & !i[1820]) | ( l_42 [7199] &  i[1820]);
assign l_41[5649]    = ( l_42 [7200] & !i[1820]) | ( l_42 [7201] &  i[1820]);
assign l_41[5650]    = ( l_42 [7202] & !i[1820]) | ( l_42 [7203] &  i[1820]);
assign l_41[5651]    = ( l_42 [7204] & !i[1820]) | ( l_42 [7205] &  i[1820]);
assign l_41[5652]    = ( l_42 [7206] & !i[1820]) | ( l_42 [7207] &  i[1820]);
assign l_41[5653]    = ( l_42 [7208] & !i[1820]) | ( l_42 [7209] &  i[1820]);
assign l_41[5654]    = ( l_42 [7210] & !i[1820]) | ( l_42 [7211] &  i[1820]);
assign l_41[5655]    = ( l_42 [7212] & !i[1820]) | ( l_42 [7213] &  i[1820]);
assign l_41[5656]    = ( l_42 [7214] & !i[1820]) | ( l_42 [7215] &  i[1820]);
assign l_41[5657]    = ( l_42 [7216] & !i[1820]) | ( l_42 [7217] &  i[1820]);
assign l_41[5658]    = ( l_42 [7218] & !i[1820]) | ( l_42 [7219] &  i[1820]);
assign l_41[5659]    = ( l_42 [7220] & !i[1820]) | ( l_42 [7221] &  i[1820]);
assign l_41[5660]    = ( l_42 [7222] & !i[1820]) | ( l_42 [7223] &  i[1820]);
assign l_41[5661]    = ( l_42 [7224] & !i[1820]) | ( l_42 [7225] &  i[1820]);
assign l_41[5662]    = ( l_42 [7226] & !i[1820]) | ( l_42 [7227] &  i[1820]);
assign l_41[5663]    = ( l_42 [7228] & !i[1820]) | ( l_42 [7229] &  i[1820]);
assign l_41[5664]    = ( l_42 [7230] & !i[1820]) | ( l_42 [7231] &  i[1820]);
assign l_41[5665]    = ( l_42 [7232] & !i[1820]) | ( l_42 [7233] &  i[1820]);
assign l_41[5666]    = ( l_42 [7234] & !i[1820]) | ( l_42 [7235] &  i[1820]);
assign l_41[5667]    = ( l_42 [7236] & !i[1820]) | ( l_42 [7237] &  i[1820]);
assign l_41[5668]    = ( l_42 [7238] & !i[1820]) | ( l_42 [7239] &  i[1820]);
assign l_41[5669]    = ( l_42 [7240] & !i[1820]) | ( l_42 [7241] &  i[1820]);
assign l_41[5670]    = ( l_42 [7242] & !i[1820]) | ( l_42 [7243] &  i[1820]);
assign l_41[5671]    = ( l_42 [7244] & !i[1820]) | ( l_42 [7245] &  i[1820]);
assign l_41[5672]    = ( l_42 [7246] & !i[1820]) | ( l_42 [7247] &  i[1820]);
assign l_41[5673]    = ( l_42 [7248] & !i[1820]) | ( l_42 [7249] &  i[1820]);
assign l_41[5674]    = ( l_42 [7250] & !i[1820]) | ( l_42 [7251] &  i[1820]);
assign l_41[5675]    = ( l_42 [7252] & !i[1820]) | ( l_42 [7253] &  i[1820]);
assign l_41[5676]    = ( l_42 [7254] & !i[1820]) | ( l_42 [7255] &  i[1820]);
assign l_41[5677]    = ( l_42 [7256] & !i[1820]) | ( l_42 [7257] &  i[1820]);
assign l_41[5678]    = ( l_42 [7258] & !i[1820]) | ( l_42 [7259] &  i[1820]);
assign l_41[5679]    = ( l_42 [7260] & !i[1820]) | ( l_42 [7261] &  i[1820]);
assign l_41[5680]    = ( l_42 [7262] & !i[1820]) | ( l_42 [7263] &  i[1820]);
assign l_41[5681]    = ( l_42 [7264] & !i[1820]) | ( l_42 [7265] &  i[1820]);
assign l_41[5682]    = ( l_42 [7266] & !i[1820]) | ( l_42 [7267] &  i[1820]);
assign l_41[5683]    = ( l_42 [7268] & !i[1820]) | ( l_42 [7269] &  i[1820]);
assign l_41[5684]    = ( l_42 [7270] & !i[1820]) | ( l_42 [7271] &  i[1820]);
assign l_41[5685]    = ( l_42 [7272] & !i[1820]) | ( l_42 [7273] &  i[1820]);
assign l_41[5686]    = ( l_42 [7274] & !i[1820]) | ( l_42 [7275] &  i[1820]);
assign l_41[5687]    = ( l_42 [7276] & !i[1820]) | ( l_42 [7277] &  i[1820]);
assign l_41[5688]    = ( l_42 [7278] & !i[1820]) | ( l_42 [7279] &  i[1820]);
assign l_41[5689]    = ( l_42 [7280] & !i[1820]) | ( l_42 [7281] &  i[1820]);
assign l_41[5690]    = ( l_42 [7282] & !i[1820]) | ( l_42 [7283] &  i[1820]);
assign l_41[5691]    = ( l_42 [7284] & !i[1820]) | ( l_42 [7285] &  i[1820]);
assign l_41[5692]    = ( l_42 [7286] & !i[1820]) | ( l_42 [7287] &  i[1820]);
assign l_41[5693]    = ( l_42 [7288] & !i[1820]) | ( l_42 [7289] &  i[1820]);
assign l_41[5694]    = ( l_42 [7290] & !i[1820]) | ( l_42 [7291] &  i[1820]);
assign l_41[5695]    = ( l_42 [7292] & !i[1820]) | ( l_42 [7293] &  i[1820]);
assign l_41[5696]    = ( l_42 [7294] & !i[1820]) | ( l_42 [7295] &  i[1820]);
assign l_41[5697]    = ( l_42 [7296] & !i[1820]) | ( l_42 [7297] &  i[1820]);
assign l_41[5698]    = ( l_42 [7298] & !i[1820]) | ( l_42 [7299] &  i[1820]);
assign l_41[5699]    = ( l_42 [7300] & !i[1820]) | ( l_42 [7301] &  i[1820]);
assign l_41[5700]    = ( l_42 [7302] & !i[1820]) | ( l_42 [7303] &  i[1820]);
assign l_41[5701]    = ( l_42 [7304] & !i[1820]) | ( l_42 [7305] &  i[1820]);
assign l_41[5702]    = ( l_42 [7306] & !i[1820]) | ( l_42 [7307] &  i[1820]);
assign l_41[5703]    = ( l_42 [7308] & !i[1820]) | ( l_42 [7309] &  i[1820]);
assign l_41[5704]    = ( l_42 [7310] & !i[1820]) | ( l_42 [7311] &  i[1820]);
assign l_41[5705]    = ( l_42 [7312] & !i[1820]) | ( l_42 [7313] &  i[1820]);
assign l_41[5706]    = ( l_42 [7314] & !i[1820]) | ( l_42 [7315] &  i[1820]);
assign l_41[5707]    = ( l_42 [7316] & !i[1820]) | ( l_42 [7317] &  i[1820]);
assign l_41[5708]    = ( l_42 [7318] & !i[1820]) | ( l_42 [7319] &  i[1820]);
assign l_41[5709]    = ( l_42 [7320] & !i[1820]) | ( l_42 [7321] &  i[1820]);
assign l_41[5710]    = ( l_42 [7322] & !i[1820]) | ( l_42 [7323] &  i[1820]);
assign l_41[5711]    = ( l_42 [7324] & !i[1820]) | ( l_42 [7325] &  i[1820]);
assign l_41[5712]    = ( l_42 [7326] & !i[1820]) | ( l_42 [7327] &  i[1820]);
assign l_41[5713]    = ( l_42 [7328] & !i[1820]) | ( l_42 [7329] &  i[1820]);
assign l_41[5714]    = ( l_42 [7330] & !i[1820]) | ( l_42 [7331] &  i[1820]);
assign l_41[5715]    = ( l_42 [7332] & !i[1820]) | ( l_42 [7333] &  i[1820]);
assign l_41[5716]    = ( l_42 [7334] & !i[1820]) | ( l_42 [7335] &  i[1820]);
assign l_41[5717]    = ( l_42 [7336] & !i[1820]) | ( l_42 [7337] &  i[1820]);
assign l_41[5718]    = ( l_42 [7338] & !i[1820]) | ( l_42 [7339] &  i[1820]);
assign l_41[5719]    = ( l_42 [7340] & !i[1820]) | ( l_42 [7341] &  i[1820]);
assign l_41[5720]    = ( l_42 [7342] & !i[1820]) | ( l_42 [7343] &  i[1820]);
assign l_41[5721]    = ( l_42 [7344] & !i[1820]) | ( l_42 [7345] &  i[1820]);
assign l_41[5722]    = ( l_42 [7346] & !i[1820]) | ( l_42 [7347] &  i[1820]);
assign l_41[5723]    = ( l_42 [7348] & !i[1820]) | ( l_42 [7349] &  i[1820]);
assign l_41[5724]    = ( l_42 [7350] & !i[1820]) | ( l_42 [7351] &  i[1820]);
assign l_41[5725]    = ( l_42 [7352] & !i[1820]) | ( l_42 [7353] &  i[1820]);
assign l_41[5726]    = ( l_42 [7354] & !i[1820]) | ( l_42 [7355] &  i[1820]);
assign l_41[5727]    = ( l_42 [7356] & !i[1820]) | ( l_42 [7357] &  i[1820]);
assign l_41[5728]    = ( l_42 [7358] & !i[1820]) | ( l_42 [7359] &  i[1820]);
assign l_41[5729]    = ( l_42 [7360] & !i[1820]) | ( l_42 [7361] &  i[1820]);
assign l_41[5730]    = ( l_42 [7362] & !i[1820]) | ( l_42 [7363] &  i[1820]);
assign l_41[5731]    = ( l_42 [7364] & !i[1820]) | ( l_42 [7365] &  i[1820]);
assign l_41[5732]    = ( l_42 [7366] & !i[1820]) | ( l_42 [7367] &  i[1820]);
assign l_41[5733]    = ( l_42 [7368] & !i[1820]) | ( l_42 [7369] &  i[1820]);
assign l_41[5734]    = ( l_42 [7370] & !i[1820]) | ( l_42 [7371] &  i[1820]);
assign l_41[5735]    = ( l_42 [7372] & !i[1820]) | ( l_42 [7373] &  i[1820]);
assign l_41[5736]    = ( l_42 [7374] & !i[1820]) | ( l_42 [7375] &  i[1820]);
assign l_41[5737]    = ( l_42 [7376] & !i[1820]) | ( l_42 [7377] &  i[1820]);
assign l_41[5738]    = ( l_42 [7378] & !i[1820]) | ( l_42 [7379] &  i[1820]);
assign l_41[5739]    = ( l_42 [7380] & !i[1820]) | ( l_42 [7381] &  i[1820]);
assign l_41[5740]    = ( l_42 [7382] & !i[1820]) | ( l_42 [7383] &  i[1820]);
assign l_41[5741]    = ( l_42 [7384] & !i[1820]) | ( l_42 [7385] &  i[1820]);
assign l_41[5742]    = ( l_42 [7386] & !i[1820]) | ( l_42 [7387] &  i[1820]);
assign l_41[5743]    = ( l_42 [7388] & !i[1820]) | ( l_42 [7389] &  i[1820]);
assign l_41[5744]    = ( l_42 [7390] & !i[1820]) | ( l_42 [7391] &  i[1820]);
assign l_41[5745]    = ( l_42 [7392] & !i[1820]) | ( l_42 [7393] &  i[1820]);
assign l_41[5746]    = ( l_42 [7394] & !i[1820]) | ( l_42 [7395] &  i[1820]);
assign l_41[5747]    = ( l_42 [7396] & !i[1820]) | ( l_42 [7397] &  i[1820]);
assign l_41[5748]    = ( l_42 [7398] & !i[1820]) | ( l_42 [7399] &  i[1820]);
assign l_41[5749]    = ( l_42 [7400] & !i[1820]) | ( l_42 [7401] &  i[1820]);
assign l_41[5750]    = ( l_42 [7402] & !i[1820]) | ( l_42 [7403] &  i[1820]);
assign l_41[5751]    = ( l_42 [7404] & !i[1820]) | ( l_42 [7405] &  i[1820]);
assign l_41[5752]    = ( l_42 [7406] & !i[1820]) | ( l_42 [7407] &  i[1820]);
assign l_41[5753]    = ( l_42 [7408] & !i[1820]) | ( l_42 [7409] &  i[1820]);
assign l_41[5754]    = ( l_42 [7410] & !i[1820]) | ( l_42 [7411] &  i[1820]);
assign l_41[5755]    = ( l_42 [7412] & !i[1820]) | ( l_42 [7413] &  i[1820]);
assign l_41[5756]    = ( l_42 [7414] & !i[1820]) | ( l_42 [7415] &  i[1820]);
assign l_41[5757]    = ( l_42 [7416] & !i[1820]) | ( l_42 [7417] &  i[1820]);
assign l_41[5758]    = ( l_42 [7418] & !i[1820]) | ( l_42 [7419] &  i[1820]);
assign l_41[5759]    = ( l_42 [7420] & !i[1820]) | ( l_42 [7421] &  i[1820]);
assign l_41[5760]    = ( l_42 [7422] & !i[1820]) | ( l_42 [7423] &  i[1820]);
assign l_41[5761]    = ( l_42 [7424] & !i[1820]) | ( l_42 [7425] &  i[1820]);
assign l_41[5762]    = ( l_42 [7426] & !i[1820]) | ( l_42 [7427] &  i[1820]);
assign l_41[5763]    = ( l_42 [7428] & !i[1820]) | ( l_42 [7429] &  i[1820]);
assign l_41[5764]    = ( l_42 [7430] & !i[1820]) | ( l_42 [7431] &  i[1820]);
assign l_41[5765]    = ( l_42 [7432] & !i[1820]) | ( l_42 [7433] &  i[1820]);
assign l_41[5766]    = ( l_42 [7434] & !i[1820]) | ( l_42 [7435] &  i[1820]);
assign l_41[5767]    = ( l_42 [7436] & !i[1820]) | ( l_42 [7437] &  i[1820]);
assign l_41[5768]    = ( l_42 [7438] & !i[1820]) | ( l_42 [7439] &  i[1820]);
assign l_41[5769]    = ( l_42 [7440] & !i[1820]) | ( l_42 [7441] &  i[1820]);
assign l_41[5770]    = ( l_42 [7442] & !i[1820]) | ( l_42 [7443] &  i[1820]);
assign l_41[5771]    = ( l_42 [7444] & !i[1820]) | ( l_42 [7445] &  i[1820]);
assign l_41[5772]    = ( l_42 [7446] & !i[1820]) | ( l_42 [7447] &  i[1820]);
assign l_41[5773]    = ( l_42 [7448] & !i[1820]) | ( l_42 [7449] &  i[1820]);
assign l_41[5774]    = ( l_42 [7450] & !i[1820]) | ( l_42 [7451] &  i[1820]);
assign l_41[5775]    = ( l_42 [7452] & !i[1820]) | ( l_42 [7453] &  i[1820]);
assign l_41[5776]    = ( l_42 [7454] & !i[1820]) | ( l_42 [7455] &  i[1820]);
assign l_41[5777]    = ( l_42 [7456] & !i[1820]) | ( l_42 [7457] &  i[1820]);
assign l_41[5778]    = ( l_42 [7458] & !i[1820]) | ( l_42 [7459] &  i[1820]);
assign l_41[5779]    = ( l_42 [7460] & !i[1820]) | ( l_42 [7461] &  i[1820]);
assign l_41[5780]    = ( l_42 [7462] & !i[1820]) | ( l_42 [7463] &  i[1820]);
assign l_41[5781]    = ( l_42 [7464] & !i[1820]) | ( l_42 [7465] &  i[1820]);
assign l_41[5782]    = ( l_42 [7466] & !i[1820]) | ( l_42 [7467] &  i[1820]);
assign l_41[5783]    = ( l_42 [7468] & !i[1820]) | ( l_42 [7469] &  i[1820]);
assign l_41[5784]    = ( l_42 [7470] & !i[1820]) | ( l_42 [7471] &  i[1820]);
assign l_41[5785]    = ( l_42 [7472] & !i[1820]) | ( l_42 [7473] &  i[1820]);
assign l_41[5786]    = ( l_42 [7474] & !i[1820]) | ( l_42 [7475] &  i[1820]);
assign l_41[5787]    = ( l_42 [7476] & !i[1820]) | ( l_42 [7477] &  i[1820]);
assign l_41[5788]    = ( l_42 [7478] & !i[1820]) | ( l_42 [7479] &  i[1820]);
assign l_41[5789]    = ( l_42 [7480] & !i[1820]) | ( l_42 [7481] &  i[1820]);
assign l_41[5790]    = ( l_42 [7482] & !i[1820]) | ( l_42 [7483] &  i[1820]);
assign l_41[5791]    = ( l_42 [7484] & !i[1820]) | ( l_42 [7485] &  i[1820]);
assign l_41[5792]    = ( l_42 [7486] & !i[1820]) | ( l_42 [7487] &  i[1820]);
assign l_41[5793]    = ( l_42 [7488] & !i[1820]) | ( l_42 [7489] &  i[1820]);
assign l_41[5794]    = ( l_42 [7490] & !i[1820]) | ( l_42 [7491] &  i[1820]);
assign l_41[5795]    = ( l_42 [7492] & !i[1820]) | ( l_42 [7493] &  i[1820]);
assign l_41[5796]    = ( l_42 [7494] & !i[1820]) | ( l_42 [7495] &  i[1820]);
assign l_41[5797]    = ( l_42 [7496] & !i[1820]) | ( l_42 [7497] &  i[1820]);
assign l_41[5798]    = ( l_42 [7498] & !i[1820]) | ( l_42 [7499] &  i[1820]);
assign l_41[5799]    = ( l_42 [7500] & !i[1820]) | ( l_42 [7501] &  i[1820]);
assign l_41[5800]    = ( l_42 [7502] & !i[1820]) | ( l_42 [7503] &  i[1820]);
assign l_41[5801]    = ( l_42 [7504] & !i[1820]) | ( l_42 [7505] &  i[1820]);
assign l_41[5802]    = ( l_42 [7506] & !i[1820]) | ( l_42 [7507] &  i[1820]);
assign l_41[5803]    = ( l_42 [7508] & !i[1820]) | ( l_42 [7509] &  i[1820]);
assign l_41[5804]    = ( l_42 [7510] & !i[1820]) | ( l_42 [7511] &  i[1820]);
assign l_41[5805]    = ( l_42 [7512] & !i[1820]) | ( l_42 [7513] &  i[1820]);
assign l_41[5806]    = ( l_42 [7514] & !i[1820]) | ( l_42 [7515] &  i[1820]);
assign l_41[5807]    = ( l_42 [7516] & !i[1820]) | ( l_42 [7517] &  i[1820]);
assign l_41[5808]    = ( l_42 [7518] & !i[1820]) | ( l_42 [7519] &  i[1820]);
assign l_41[5809]    = ( l_42 [7520] & !i[1820]) | ( l_42 [7521] &  i[1820]);
assign l_41[5810]    = ( l_42 [7522] & !i[1820]) | ( l_42 [7523] &  i[1820]);
assign l_41[5811]    = ( l_42 [7524] & !i[1820]) | ( l_42 [7525] &  i[1820]);
assign l_41[5812]    = ( l_42 [7526] & !i[1820]) | ( l_42 [7527] &  i[1820]);
assign l_41[5813]    = ( l_42 [7528] & !i[1820]) | ( l_42 [7529] &  i[1820]);
assign l_41[5814]    = ( l_42 [7530] & !i[1820]) | ( l_42 [7531] &  i[1820]);
assign l_41[5815]    = ( l_42 [7532] & !i[1820]) | ( l_42 [7533] &  i[1820]);
assign l_41[5816]    = ( l_42 [7534] & !i[1820]) | ( l_42 [7535] &  i[1820]);
assign l_41[5817]    = ( l_42 [7536] & !i[1820]) | ( l_42 [7537] &  i[1820]);
assign l_41[5818]    = ( l_42 [7538] & !i[1820]) | ( l_42 [7539] &  i[1820]);
assign l_41[5819]    = ( l_42 [7540] & !i[1820]) | ( l_42 [7541] &  i[1820]);
assign l_41[5820]    = ( l_42 [7542] & !i[1820]) | ( l_42 [7543] &  i[1820]);
assign l_41[5821]    = ( l_42 [7544] & !i[1820]) | ( l_42 [7545] &  i[1820]);
assign l_41[5822]    = ( l_42 [7546] & !i[1820]) | ( l_42 [7547] &  i[1820]);
assign l_41[5823]    = ( l_42 [7548] & !i[1820]) | ( l_42 [7549] &  i[1820]);
assign l_41[5824]    = ( l_42 [7550] & !i[1820]) | ( l_42 [7551] &  i[1820]);
assign l_41[5825]    = ( l_42 [7552] & !i[1820]) | ( l_42 [7553] &  i[1820]);
assign l_41[5826]    = ( l_42 [7554] & !i[1820]) | ( l_42 [7555] &  i[1820]);
assign l_41[5827]    = ( l_42 [7556] & !i[1820]) | ( l_42 [7557] &  i[1820]);
assign l_41[5828]    = ( l_42 [7558] & !i[1820]) | ( l_42 [7559] &  i[1820]);
assign l_41[5829]    = ( l_42 [7560] & !i[1820]) | ( l_42 [7561] &  i[1820]);
assign l_41[5830]    = ( l_42 [7562] & !i[1820]) | ( l_42 [7563] &  i[1820]);
assign l_41[5831]    = ( l_42 [7564] & !i[1820]) | ( l_42 [7565] &  i[1820]);
assign l_41[5832]    = ( l_42 [7566] & !i[1820]) | ( l_42 [7567] &  i[1820]);
assign l_41[5833]    = ( l_42 [7568] & !i[1820]) | ( l_42 [7569] &  i[1820]);
assign l_41[5834]    = ( l_42 [7570] & !i[1820]) | ( l_42 [7571] &  i[1820]);
assign l_41[5835]    = ( l_42 [7572] & !i[1820]) | ( l_42 [7573] &  i[1820]);
assign l_41[5836]    = ( l_42 [7574] & !i[1820]) | ( l_42 [7575] &  i[1820]);
assign l_41[5837]    = ( l_42 [7576] & !i[1820]) | ( l_42 [7577] &  i[1820]);
assign l_41[5838]    = ( l_42 [7578] & !i[1820]) | ( l_42 [7579] &  i[1820]);
assign l_41[5839]    = ( l_42 [7580] & !i[1820]) | ( l_42 [7581] &  i[1820]);
assign l_41[5840]    = ( l_42 [7582] & !i[1820]) | ( l_42 [7583] &  i[1820]);
assign l_41[5841]    = ( l_42 [7584] & !i[1820]) | ( l_42 [7585] &  i[1820]);
assign l_41[5842]    = ( l_42 [7586] & !i[1820]) | ( l_42 [7587] &  i[1820]);
assign l_41[5843]    = ( l_42 [7588] & !i[1820]) | ( l_42 [7589] &  i[1820]);
assign l_41[5844]    = ( l_42 [7590] & !i[1820]) | ( l_42 [7591] &  i[1820]);
assign l_41[5845]    = ( l_42 [7592] & !i[1820]) | ( l_42 [7593] &  i[1820]);
assign l_41[5846]    = ( l_42 [7594] & !i[1820]) | ( l_42 [7595] &  i[1820]);
assign l_41[5847]    = ( l_42 [7596] & !i[1820]) | ( l_42 [7597] &  i[1820]);
assign l_41[5848]    = ( l_42 [7598] & !i[1820]) | ( l_42 [7599] &  i[1820]);
assign l_41[5849]    = ( l_42 [7600] & !i[1820]) | ( l_42 [7601] &  i[1820]);
assign l_41[5850]    = ( l_42 [7602] & !i[1820]) | ( l_42 [7603] &  i[1820]);
assign l_41[5851]    = ( l_42 [7604] & !i[1820]) | ( l_42 [7605] &  i[1820]);
assign l_41[5852]    = ( l_42 [7606] & !i[1820]) | ( l_42 [7607] &  i[1820]);
assign l_41[5853]    = ( l_42 [7608] & !i[1820]) | ( l_42 [7609] &  i[1820]);
assign l_41[5854]    = ( l_42 [7610] & !i[1820]) | ( l_42 [7611] &  i[1820]);
assign l_41[5855]    = ( l_42 [7612] & !i[1820]) | ( l_42 [7613] &  i[1820]);
assign l_41[5856]    = ( l_42 [7614] & !i[1820]) | ( l_42 [7615] &  i[1820]);
assign l_41[5857]    = ( l_42 [7616] & !i[1820]) | ( l_42 [7617] &  i[1820]);
assign l_41[5858]    = ( l_42 [7618] & !i[1820]) | ( l_42 [7619] &  i[1820]);
assign l_41[5859]    = ( l_42 [7620] & !i[1820]) | ( l_42 [7621] &  i[1820]);
assign l_41[5860]    = ( l_42 [7622] & !i[1820]) | ( l_42 [7623] &  i[1820]);
assign l_41[5861]    = ( l_42 [7624] & !i[1820]) | ( l_42 [7625] &  i[1820]);
assign l_41[5862]    = ( l_42 [7626] & !i[1820]) | ( l_42 [7627] &  i[1820]);
assign l_41[5863]    = ( l_42 [7628] & !i[1820]) | ( l_42 [7629] &  i[1820]);
assign l_41[5864]    = ( l_42 [7630] & !i[1820]) | ( l_42 [7631] &  i[1820]);
assign l_41[5865]    = ( l_42 [7632] & !i[1820]) | ( l_42 [7633] &  i[1820]);
assign l_41[5866]    = ( l_42 [7634] & !i[1820]) | ( l_42 [7635] &  i[1820]);
assign l_41[5867]    = ( l_42 [7636] & !i[1820]) | ( l_42 [7637] &  i[1820]);
assign l_41[5868]    = ( l_42 [7638] & !i[1820]) | ( l_42 [7639] &  i[1820]);
assign l_41[5869]    = ( l_42 [7640] & !i[1820]) | ( l_42 [7641] &  i[1820]);
assign l_41[5870]    = ( l_42 [7642] & !i[1820]) | ( l_42 [7643] &  i[1820]);
assign l_41[5871]    = ( l_42 [7644] & !i[1820]) | ( l_42 [7645] &  i[1820]);
assign l_41[5872]    = ( l_42 [7646] & !i[1820]) | ( l_42 [7647] &  i[1820]);
assign l_41[5873]    = ( l_42 [7648] & !i[1820]) | ( l_42 [7649] &  i[1820]);
assign l_41[5874]    = ( l_42 [7650] & !i[1820]) | ( l_42 [7651] &  i[1820]);
assign l_41[5875]    = ( l_42 [7652] & !i[1820]) | ( l_42 [7653] &  i[1820]);
assign l_41[5876]    = ( l_42 [7654] & !i[1820]) | ( l_42 [7655] &  i[1820]);
assign l_41[5877]    = ( l_42 [7656] & !i[1820]) | ( l_42 [7657] &  i[1820]);
assign l_41[5878]    = ( l_42 [7658] & !i[1820]) | ( l_42 [7659] &  i[1820]);
assign l_41[5879]    = ( l_42 [7660] & !i[1820]) | ( l_42 [7661] &  i[1820]);
assign l_41[5880]    = ( l_42 [7662] & !i[1820]) | ( l_42 [7663] &  i[1820]);
assign l_41[5881]    = ( l_42 [7664] & !i[1820]) | ( l_42 [7665] &  i[1820]);
assign l_41[5882]    = ( l_42 [7666] & !i[1820]) | ( l_42 [7667] &  i[1820]);
assign l_41[5883]    = ( l_42 [7668] & !i[1820]) | ( l_42 [7669] &  i[1820]);
assign l_41[5884]    = ( l_42 [7670] & !i[1820]) | ( l_42 [7671] &  i[1820]);
assign l_41[5885]    = ( l_42 [7672] & !i[1820]) | ( l_42 [7673] &  i[1820]);
assign l_41[5886]    = ( l_42 [7674] & !i[1820]) | ( l_42 [7675] &  i[1820]);
assign l_41[5887]    = ( l_42 [7676] & !i[1820]) | ( l_42 [7677] &  i[1820]);
assign l_41[5888]    = ( l_42 [7678] & !i[1820]) | ( l_42 [7679] &  i[1820]);
assign l_41[5889]    = ( l_42 [7680] & !i[1820]) | ( l_42 [7681] &  i[1820]);
assign l_41[5890]    = ( l_42 [7682] & !i[1820]) | ( l_42 [7683] &  i[1820]);
assign l_41[5891]    = ( l_42 [7684] & !i[1820]) | ( l_42 [7685] &  i[1820]);
assign l_41[5892]    = ( l_42 [7686] & !i[1820]) | ( l_42 [7687] &  i[1820]);
assign l_41[5893]    = ( l_42 [7688] & !i[1820]) | ( l_42 [7689] &  i[1820]);
assign l_41[5894]    = ( l_42 [7690] & !i[1820]) | ( l_42 [7691] &  i[1820]);
assign l_41[5895]    = ( l_42 [7692] & !i[1820]) | ( l_42 [7693] &  i[1820]);
assign l_41[5896]    = ( l_42 [7694] & !i[1820]) | ( l_42 [7695] &  i[1820]);
assign l_41[5897]    = ( l_42 [7696] & !i[1820]) | ( l_42 [7697] &  i[1820]);
assign l_41[5898]    = ( l_42 [7698] & !i[1820]) | ( l_42 [7699] &  i[1820]);
assign l_41[5899]    = ( l_42 [7700] & !i[1820]) | ( l_42 [7701] &  i[1820]);
assign l_41[5900]    = ( l_42 [7702] & !i[1820]) | ( l_42 [7703] &  i[1820]);
assign l_41[5901]    = ( l_42 [7704] & !i[1820]) | ( l_42 [7705] &  i[1820]);
assign l_41[5902]    = ( l_42 [7706] & !i[1820]) | ( l_42 [7707] &  i[1820]);
assign l_41[5903]    = ( l_42 [7708] & !i[1820]) | ( l_42 [7709] &  i[1820]);
assign l_41[5904]    = ( l_42 [7710] & !i[1820]) | ( l_42 [7711] &  i[1820]);
assign l_41[5905]    = ( l_42 [7712] & !i[1820]) | ( l_42 [7713] &  i[1820]);
assign l_41[5906]    = ( l_42 [7714] & !i[1820]) | ( l_42 [7715] &  i[1820]);
assign l_41[5907]    = ( l_42 [7716] & !i[1820]) | ( l_42 [7717] &  i[1820]);
assign l_41[5908]    = ( l_42 [7718] & !i[1820]) | ( l_42 [7719] &  i[1820]);
assign l_41[5909]    = ( l_42 [7720] & !i[1820]) | ( l_42 [7721] &  i[1820]);
assign l_41[5910]    = ( l_42 [7722] & !i[1820]) | ( l_42 [7723] &  i[1820]);
assign l_41[5911]    = ( l_42 [7724] & !i[1820]) | ( l_42 [7725] &  i[1820]);
assign l_41[5912]    = ( l_42 [7726] & !i[1820]) | ( l_42 [7727] &  i[1820]);
assign l_41[5913]    = ( l_42 [7728] & !i[1820]) | ( l_42 [7729] &  i[1820]);
assign l_41[5914]    = ( l_42 [7730] & !i[1820]) | ( l_42 [7731] &  i[1820]);
assign l_41[5915]    = ( l_42 [7732] & !i[1820]) | ( l_42 [7733] &  i[1820]);
assign l_41[5916]    = ( l_42 [7734] & !i[1820]) | ( l_42 [7735] &  i[1820]);
assign l_41[5917]    = ( l_42 [7736] & !i[1820]) | ( l_42 [7737] &  i[1820]);
assign l_41[5918]    = ( l_42 [7738] & !i[1820]) | ( l_42 [7739] &  i[1820]);
assign l_41[5919]    = ( l_42 [7740] & !i[1820]) | ( l_42 [7741] &  i[1820]);
assign l_41[5920]    = ( l_42 [7742] & !i[1820]) | ( l_42 [7743] &  i[1820]);
assign l_41[5921]    = ( l_42 [7744] & !i[1820]) | ( l_42 [7745] &  i[1820]);
assign l_41[5922]    = ( l_42 [7746] & !i[1820]) | ( l_42 [7747] &  i[1820]);
assign l_41[5923]    = ( l_42 [7748] & !i[1820]) | ( l_42 [7749] &  i[1820]);
assign l_41[5924]    = ( l_42 [7750] & !i[1820]) | ( l_42 [7751] &  i[1820]);
assign l_41[5925]    = ( l_42 [7752] & !i[1820]) | ( l_42 [7753] &  i[1820]);
assign l_41[5926]    = ( l_42 [7754] & !i[1820]) | ( l_42 [7755] &  i[1820]);
assign l_41[5927]    = ( l_42 [7756] & !i[1820]) | ( l_42 [7757] &  i[1820]);
assign l_41[5928]    = ( l_42 [7758] & !i[1820]) | ( l_42 [7759] &  i[1820]);
assign l_41[5929]    = ( l_42 [7760] & !i[1820]) | ( l_42 [7761] &  i[1820]);
assign l_41[5930]    = ( l_42 [7762] & !i[1820]) | ( l_42 [7763] &  i[1820]);
assign l_41[5931]    = ( l_42 [7764] & !i[1820]) | ( l_42 [7765] &  i[1820]);
assign l_41[5932]    = ( l_42 [7766] & !i[1820]) | ( l_42 [7767] &  i[1820]);
assign l_41[5933]    = ( l_42 [7768] & !i[1820]) | ( l_42 [7769] &  i[1820]);
assign l_41[5934]    = ( l_42 [7770] & !i[1820]) | ( l_42 [7771] &  i[1820]);
assign l_41[5935]    = ( l_42 [7772] & !i[1820]) | ( l_42 [7773] &  i[1820]);
assign l_41[5936]    = ( l_42 [7774] & !i[1820]) | ( l_42 [7775] &  i[1820]);
assign l_41[5937]    = ( l_42 [7776] & !i[1820]) | ( l_42 [7777] &  i[1820]);
assign l_41[5938]    = ( l_42 [7778] & !i[1820]) | ( l_42 [7779] &  i[1820]);
assign l_41[5939]    = ( l_42 [7780] & !i[1820]) | ( l_42 [7781] &  i[1820]);
assign l_41[5940]    = ( l_42 [7782] & !i[1820]) | ( l_42 [7783] &  i[1820]);
assign l_41[5941]    = ( l_42 [7784] & !i[1820]) | ( l_42 [7785] &  i[1820]);
assign l_41[5942]    = ( l_42 [7786] & !i[1820]) | ( l_42 [7787] &  i[1820]);
assign l_41[5943]    = ( l_42 [7788] & !i[1820]) | ( l_42 [7789] &  i[1820]);
assign l_41[5944]    = ( l_42 [7790] & !i[1820]) | ( l_42 [7791] &  i[1820]);
assign l_41[5945]    = ( l_42 [7792] & !i[1820]) | ( l_42 [7793] &  i[1820]);
assign l_41[5946]    = ( l_42 [7794] & !i[1820]) | ( l_42 [7795] &  i[1820]);
assign l_41[5947]    = ( l_42 [7796] & !i[1820]) | ( l_42 [7797] &  i[1820]);
assign l_41[5948]    = ( l_42 [7798] & !i[1820]) | ( l_42 [7799] &  i[1820]);
assign l_41[5949]    = ( l_42 [7800] & !i[1820]) | ( l_42 [7801] &  i[1820]);
assign l_41[5950]    = ( l_42 [7802] & !i[1820]) | ( l_42 [7803] &  i[1820]);
assign l_41[5951]    = ( l_42 [7804] & !i[1820]) | ( l_42 [7805] &  i[1820]);
assign l_41[5952]    = ( l_42 [7806] & !i[1820]) | ( l_42 [7807] &  i[1820]);
assign l_41[5953]    = ( l_42 [7808] & !i[1820]) | ( l_42 [7809] &  i[1820]);
assign l_41[5954]    = ( l_42 [7810] & !i[1820]) | ( l_42 [7811] &  i[1820]);
assign l_41[5955]    = ( l_42 [7812] & !i[1820]) | ( l_42 [7813] &  i[1820]);
assign l_41[5956]    = ( l_42 [7814] & !i[1820]) | ( l_42 [7815] &  i[1820]);
assign l_41[5957]    = ( l_42 [7816] & !i[1820]) | ( l_42 [7817] &  i[1820]);
assign l_41[5958]    = ( l_42 [7818] & !i[1820]) | ( l_42 [7819] &  i[1820]);
assign l_41[5959]    = ( l_42 [7820] & !i[1820]) | ( l_42 [7821] &  i[1820]);
assign l_41[5960]    = ( l_42 [7822] & !i[1820]) | ( l_42 [7823] &  i[1820]);
assign l_41[5961]    = ( l_42 [7824] & !i[1820]) | ( l_42 [7825] &  i[1820]);
assign l_41[5962]    = ( l_42 [7826] & !i[1820]) | ( l_42 [7827] &  i[1820]);
assign l_41[5963]    = ( l_42 [7828] & !i[1820]) | ( l_42 [7829] &  i[1820]);
assign l_41[5964]    = ( l_42 [7830] & !i[1820]) | ( l_42 [7831] &  i[1820]);
assign l_41[5965]    = ( l_42 [7832] & !i[1820]) | ( l_42 [7833] &  i[1820]);
assign l_41[5966]    = ( l_42 [7834] & !i[1820]) | ( l_42 [7835] &  i[1820]);
assign l_41[5967]    = ( l_42 [7836] & !i[1820]) | ( l_42 [7837] &  i[1820]);
assign l_41[5968]    = ( l_42 [7838] & !i[1820]) | ( l_42 [7839] &  i[1820]);
assign l_41[5969]    = ( l_42 [7840] & !i[1820]) | ( l_42 [7841] &  i[1820]);
assign l_41[5970]    = ( l_42 [7842] & !i[1820]) | ( l_42 [7843] &  i[1820]);
assign l_41[5971]    = ( l_42 [7844] & !i[1820]) | ( l_42 [7845] &  i[1820]);
assign l_41[5972]    = ( l_42 [7846] & !i[1820]) | ( l_42 [7847] &  i[1820]);
assign l_41[5973]    = ( l_42 [7848] & !i[1820]) | ( l_42 [7849] &  i[1820]);
assign l_41[5974]    = ( l_42 [7850] & !i[1820]) | ( l_42 [7851] &  i[1820]);
assign l_41[5975]    = ( l_42 [7852] & !i[1820]) | ( l_42 [7853] &  i[1820]);
assign l_41[5976]    = ( l_42 [7854] & !i[1820]) | ( l_42 [7855] &  i[1820]);
assign l_41[5977]    = ( l_42 [7856] & !i[1820]) | ( l_42 [7857] &  i[1820]);
assign l_41[5978]    = ( l_42 [7858] & !i[1820]) | ( l_42 [7859] &  i[1820]);
assign l_41[5979]    = ( l_42 [7860] & !i[1820]) | ( l_42 [7861] &  i[1820]);
assign l_41[5980]    = ( l_42 [7862] & !i[1820]) | ( l_42 [7863] &  i[1820]);
assign l_41[5981]    = ( l_42 [7864] & !i[1820]) | ( l_42 [7865] &  i[1820]);
assign l_41[5982]    = ( l_42 [7866] & !i[1820]) | ( l_42 [7867] &  i[1820]);
assign l_41[5983]    = ( l_42 [7868] & !i[1820]) | ( l_42 [7869] &  i[1820]);
assign l_41[5984]    = ( l_42 [7870] & !i[1820]) | ( l_42 [7871] &  i[1820]);
assign l_41[5985]    = ( l_42 [7872] & !i[1820]) | ( l_42 [7873] &  i[1820]);
assign l_41[5986]    = ( l_42 [7874] & !i[1820]) | ( l_42 [7875] &  i[1820]);
assign l_41[5987]    = ( l_42 [7876] & !i[1820]) | ( l_42 [7877] &  i[1820]);
assign l_41[5988]    = ( l_42 [7878] & !i[1820]) | ( l_42 [7879] &  i[1820]);
assign l_41[5989]    = ( l_42 [7880] & !i[1820]) | ( l_42 [7881] &  i[1820]);
assign l_41[5990]    = ( l_42 [7882] & !i[1820]) | ( l_42 [7883] &  i[1820]);
assign l_41[5991]    = ( l_42 [7884] & !i[1820]) | ( l_42 [7885] &  i[1820]);
assign l_41[5992]    = ( l_42 [7886] & !i[1820]) | ( l_42 [7887] &  i[1820]);
assign l_41[5993]    = ( l_42 [7888] & !i[1820]) | ( l_42 [7889] &  i[1820]);
assign l_41[5994]    = ( l_42 [7890] & !i[1820]) | ( l_42 [7891] &  i[1820]);
assign l_41[5995]    = ( l_42 [7892] & !i[1820]) | ( l_42 [7893] &  i[1820]);
assign l_41[5996]    = ( l_42 [7894] & !i[1820]) | ( l_42 [7895] &  i[1820]);
assign l_41[5997]    = ( l_42 [7896] & !i[1820]) | ( l_42 [7897] &  i[1820]);
assign l_41[5998]    = ( l_42 [7898] & !i[1820]) | ( l_42 [7899] &  i[1820]);
assign l_41[5999]    = ( l_42 [7900] & !i[1820]) | ( l_42 [7901] &  i[1820]);
assign l_41[6000]    = ( l_42 [7902] & !i[1820]) | ( l_42 [7903] &  i[1820]);
assign l_41[6001]    = ( l_42 [7904] & !i[1820]) | ( l_42 [7905] &  i[1820]);
assign l_41[6002]    = ( l_42 [7906] & !i[1820]) | ( l_42 [7907] &  i[1820]);
assign l_41[6003]    = ( l_42 [7908] & !i[1820]) | ( l_42 [7909] &  i[1820]);
assign l_41[6004]    = ( l_42 [7910] & !i[1820]) | ( l_42 [7911] &  i[1820]);
assign l_41[6005]    = ( l_42 [7912] & !i[1820]) | ( l_42 [7913] &  i[1820]);
assign l_41[6006]    = ( l_42 [7914] & !i[1820]) | ( l_42 [7915] &  i[1820]);
assign l_41[6007]    = ( l_42 [7916] & !i[1820]) | ( l_42 [7917] &  i[1820]);
assign l_41[6008]    = ( l_42 [7918] & !i[1820]) | ( l_42 [7919] &  i[1820]);
assign l_41[6009]    = ( l_42 [7920] & !i[1820]) | ( l_42 [7921] &  i[1820]);
assign l_41[6010]    = ( l_42 [7922] & !i[1820]) | ( l_42 [7923] &  i[1820]);
assign l_41[6011]    = ( l_42 [7924] & !i[1820]) | ( l_42 [7925] &  i[1820]);
assign l_41[6012]    = ( l_42 [7926] & !i[1820]) | ( l_42 [7927] &  i[1820]);
assign l_41[6013]    = ( l_42 [7928] & !i[1820]) | ( l_42 [7929] &  i[1820]);
assign l_41[6014]    = ( l_42 [7930] & !i[1820]) | ( l_42 [7931] &  i[1820]);
assign l_41[6015]    = ( l_42 [7932] & !i[1820]) | ( l_42 [7933] &  i[1820]);
assign l_41[6016]    = ( l_42 [7934] & !i[1820]) | ( l_42 [7935] &  i[1820]);
assign l_41[6017]    = ( l_42 [7936] & !i[1820]) | ( l_42 [7937] &  i[1820]);
assign l_41[6018]    = ( l_42 [7938] & !i[1820]) | ( l_42 [7939] &  i[1820]);
assign l_41[6019]    = ( l_42 [7940] & !i[1820]) | ( l_42 [7941] &  i[1820]);
assign l_41[6020]    = ( l_42 [7942] & !i[1820]) | ( l_42 [7943] &  i[1820]);
assign l_41[6021]    = ( l_42 [7944] & !i[1820]) | ( l_42 [7945] &  i[1820]);
assign l_41[6022]    = ( l_42 [7946] & !i[1820]) | ( l_42 [7947] &  i[1820]);
assign l_41[6023]    = ( l_42 [7948] & !i[1820]) | ( l_42 [7949] &  i[1820]);
assign l_41[6024]    = ( l_42 [7950] & !i[1820]) | ( l_42 [7951] &  i[1820]);
assign l_41[6025]    = ( l_42 [7952] & !i[1820]) | ( l_42 [7953] &  i[1820]);
assign l_41[6026]    = ( l_42 [7954] & !i[1820]) | ( l_42 [7955] &  i[1820]);
assign l_41[6027]    = ( l_42 [7956] & !i[1820]) | ( l_42 [7957] &  i[1820]);
assign l_41[6028]    = ( l_42 [7958] & !i[1820]) | ( l_42 [7959] &  i[1820]);
assign l_41[6029]    = ( l_42 [7960] & !i[1820]) | ( l_42 [7961] &  i[1820]);
assign l_41[6030]    = ( l_42 [7962] & !i[1820]) | ( l_42 [7963] &  i[1820]);
assign l_41[6031]    = ( l_42 [7964] & !i[1820]) | ( l_42 [7965] &  i[1820]);
assign l_41[6032]    = ( l_42 [7966] & !i[1820]) | ( l_42 [7967] &  i[1820]);
assign l_41[6033]    = ( l_42 [7968] & !i[1820]) | ( l_42 [7969] &  i[1820]);
assign l_41[6034]    = ( l_42 [7970] & !i[1820]) | ( l_42 [7971] &  i[1820]);
assign l_41[6035]    = ( l_42 [7972] & !i[1820]) | ( l_42 [7973] &  i[1820]);
assign l_41[6036]    = ( l_42 [7974] & !i[1820]) | ( l_42 [7975] &  i[1820]);
assign l_41[6037]    = ( l_42 [7976] & !i[1820]) | ( l_42 [7977] &  i[1820]);
assign l_41[6038]    = ( l_42 [7978] & !i[1820]) | ( l_42 [7979] &  i[1820]);
assign l_41[6039]    = ( l_42 [7980] & !i[1820]) | ( l_42 [7981] &  i[1820]);
assign l_41[6040]    = ( l_42 [7982] & !i[1820]) | ( l_42 [7983] &  i[1820]);
assign l_41[6041]    = ( l_42 [7984] & !i[1820]) | ( l_42 [7985] &  i[1820]);
assign l_41[6042]    = ( l_42 [7986] & !i[1820]) | ( l_42 [7987] &  i[1820]);
assign l_41[6043]    = ( l_42 [7988] & !i[1820]) | ( l_42 [7989] &  i[1820]);
assign l_41[6044]    = ( l_42 [7990] & !i[1820]) | ( l_42 [7991] &  i[1820]);
assign l_41[6045]    = ( l_42 [7992] & !i[1820]) | ( l_42 [7993] &  i[1820]);
assign l_41[6046]    = ( l_42 [7994] & !i[1820]) | ( l_42 [7995] &  i[1820]);
assign l_41[6047]    = ( l_42 [7996] & !i[1820]) | ( l_42 [7997] &  i[1820]);
assign l_41[6048]    = ( l_42 [7998] & !i[1820]) | ( l_42 [7999] &  i[1820]);
assign l_41[6049]    = ( l_42 [8000] & !i[1820]) | ( l_42 [8001] &  i[1820]);
assign l_41[6050]    = ( l_42 [8002] & !i[1820]) | ( l_42 [8003] &  i[1820]);
assign l_41[6051]    = ( l_42 [8004] & !i[1820]) | ( l_42 [8005] &  i[1820]);
assign l_41[6052]    = ( l_42 [8006] & !i[1820]) | ( l_42 [8007] &  i[1820]);
assign l_41[6053]    = ( l_42 [8008] & !i[1820]) | ( l_42 [8009] &  i[1820]);
assign l_41[6054]    = ( l_42 [8010] & !i[1820]) | ( l_42 [8011] &  i[1820]);
assign l_41[6055]    = ( l_42 [8012] & !i[1820]) | ( l_42 [8013] &  i[1820]);
assign l_41[6056]    = ( l_42 [8014] & !i[1820]) | ( l_42 [8015] &  i[1820]);
assign l_41[6057]    = ( l_42 [8016] & !i[1820]) | ( l_42 [8017] &  i[1820]);
assign l_41[6058]    = ( l_42 [8018] & !i[1820]) | ( l_42 [8019] &  i[1820]);
assign l_41[6059]    = ( l_42 [8020] & !i[1820]) | ( l_42 [8021] &  i[1820]);
assign l_41[6060]    = ( l_42 [8022] & !i[1820]) | ( l_42 [8023] &  i[1820]);
assign l_41[6061]    = ( l_42 [8024] & !i[1820]) | ( l_42 [8025] &  i[1820]);
assign l_41[6062]    = ( l_42 [8026] & !i[1820]) | ( l_42 [8027] &  i[1820]);
assign l_41[6063]    = ( l_42 [8028] & !i[1820]) | ( l_42 [8029] &  i[1820]);
assign l_41[6064]    = ( l_42 [8030] & !i[1820]) | ( l_42 [8031] &  i[1820]);
assign l_41[6065]    = ( l_42 [8032] & !i[1820]) | ( l_42 [8033] &  i[1820]);
assign l_41[6066]    = ( l_42 [8034] & !i[1820]) | ( l_42 [8035] &  i[1820]);
assign l_41[6067]    = ( l_42 [8036] & !i[1820]) | ( l_42 [8037] &  i[1820]);
assign l_41[6068]    = ( l_42 [8038] & !i[1820]) | ( l_42 [8039] &  i[1820]);
assign l_41[6069]    = ( l_42 [8040] & !i[1820]) | ( l_42 [8041] &  i[1820]);
assign l_41[6070]    = ( l_42 [8042] & !i[1820]) | ( l_42 [8043] &  i[1820]);
assign l_41[6071]    = ( l_42 [8044] & !i[1820]) | ( l_42 [8045] &  i[1820]);
assign l_41[6072]    = ( l_42 [8046] & !i[1820]) | ( l_42 [8047] &  i[1820]);
assign l_41[6073]    = ( l_42 [8048] & !i[1820]) | ( l_42 [8049] &  i[1820]);
assign l_41[6074]    = ( l_42 [8050] & !i[1820]) | ( l_42 [8051] &  i[1820]);
assign l_41[6075]    = ( l_42 [8052] & !i[1820]) | ( l_42 [8053] &  i[1820]);
assign l_41[6076]    = ( l_42 [8054] & !i[1820]) | ( l_42 [8055] &  i[1820]);
assign l_41[6077]    = ( l_42 [8056] & !i[1820]) | ( l_42 [8057] &  i[1820]);
assign l_41[6078]    = ( l_42 [8058] & !i[1820]) | ( l_42 [8059] &  i[1820]);
assign l_41[6079]    = ( l_42 [8060] & !i[1820]) | ( l_42 [8061] &  i[1820]);
assign l_41[6080]    = ( l_42 [8062] & !i[1820]) | ( l_42 [8063] &  i[1820]);
assign l_41[6081]    = ( l_42 [8064] & !i[1820]) | ( l_42 [8065] &  i[1820]);
assign l_41[6082]    = ( l_42 [8066] & !i[1820]) | ( l_42 [8067] &  i[1820]);
assign l_41[6083]    = ( l_42 [8068] & !i[1820]) | ( l_42 [8069] &  i[1820]);
assign l_41[6084]    = ( l_42 [8070] & !i[1820]) | ( l_42 [8071] &  i[1820]);
assign l_41[6085]    = ( l_42 [8072] & !i[1820]) | ( l_42 [8073] &  i[1820]);
assign l_41[6086]    = ( l_42 [8074] & !i[1820]) | ( l_42 [8075] &  i[1820]);
assign l_41[6087]    = ( l_42 [8076] & !i[1820]) | ( l_42 [8077] &  i[1820]);
assign l_41[6088]    = ( l_42 [8078] & !i[1820]) | ( l_42 [8079] &  i[1820]);
assign l_41[6089]    = ( l_42 [8080] & !i[1820]) | ( l_42 [8081] &  i[1820]);
assign l_41[6090]    = ( l_42 [8082] & !i[1820]) | ( l_42 [8083] &  i[1820]);
assign l_41[6091]    = ( l_42 [8084] & !i[1820]) | ( l_42 [8085] &  i[1820]);
assign l_41[6092]    = ( l_42 [8086] & !i[1820]) | ( l_42 [8087] &  i[1820]);
assign l_41[6093]    = ( l_42 [8088] & !i[1820]) | ( l_42 [8089] &  i[1820]);
assign l_41[6094]    = ( l_42 [8090] & !i[1820]) | ( l_42 [8091] &  i[1820]);
assign l_41[6095]    = ( l_42 [8092] & !i[1820]) | ( l_42 [8093] &  i[1820]);
assign l_41[6096]    = ( l_42 [8094] & !i[1820]) | ( l_42 [8095] &  i[1820]);
assign l_41[6097]    = ( l_42 [8096] & !i[1820]) | ( l_42 [8097] &  i[1820]);
assign l_41[6098]    = ( l_42 [8098] & !i[1820]) | ( l_42 [8099] &  i[1820]);
assign l_41[6099]    = ( l_42 [8100] & !i[1820]) | ( l_42 [8101] &  i[1820]);
assign l_41[6100]    = ( l_42 [8102] & !i[1820]) | ( l_42 [8103] &  i[1820]);
assign l_41[6101]    = ( l_42 [8104] & !i[1820]) | ( l_42 [8105] &  i[1820]);
assign l_41[6102]    = ( l_42 [8106] & !i[1820]) | ( l_42 [8107] &  i[1820]);
assign l_41[6103]    = ( l_42 [8108] & !i[1820]) | ( l_42 [8109] &  i[1820]);
assign l_41[6104]    = ( l_42 [8110] & !i[1820]) | ( l_42 [8111] &  i[1820]);
assign l_41[6105]    = ( l_42 [8112] & !i[1820]) | ( l_42 [8113] &  i[1820]);
assign l_41[6106]    = ( l_42 [8114] & !i[1820]) | ( l_42 [8115] &  i[1820]);
assign l_41[6107]    = ( l_42 [8116] & !i[1820]) | ( l_42 [8117] &  i[1820]);
assign l_41[6108]    = ( l_42 [8118] & !i[1820]) | ( l_42 [8119] &  i[1820]);
assign l_41[6109]    = ( l_42 [8120] & !i[1820]) | ( l_42 [8121] &  i[1820]);
assign l_41[6110]    = ( l_42 [8122] & !i[1820]) | ( l_42 [8123] &  i[1820]);
assign l_41[6111]    = ( l_42 [8124] & !i[1820]) | ( l_42 [8125] &  i[1820]);
assign l_41[6112]    = ( l_42 [8126] & !i[1820]) | ( l_42 [8127] &  i[1820]);
assign l_41[6113]    = ( l_42 [8128] & !i[1820]) | ( l_42 [8129] &  i[1820]);
assign l_41[6114]    = ( l_42 [8130] & !i[1820]) | ( l_42 [8131] &  i[1820]);
assign l_41[6115]    = ( l_42 [8132] & !i[1820]) | ( l_42 [8133] &  i[1820]);
assign l_41[6116]    = ( l_42 [8134] & !i[1820]) | ( l_42 [8135] &  i[1820]);
assign l_41[6117]    = ( l_42 [8136] & !i[1820]) | ( l_42 [8137] &  i[1820]);
assign l_41[6118]    = ( l_42 [8138] & !i[1820]) | ( l_42 [8139] &  i[1820]);
assign l_41[6119]    = ( l_42 [8140] & !i[1820]) | ( l_42 [8141] &  i[1820]);
assign l_41[6120]    = ( l_42 [8142] & !i[1820]) | ( l_42 [8143] &  i[1820]);
assign l_41[6121]    = ( l_42 [8144] & !i[1820]) | ( l_42 [8145] &  i[1820]);
assign l_41[6122]    = ( l_42 [8146] & !i[1820]) | ( l_42 [8147] &  i[1820]);
assign l_41[6123]    = ( l_42 [8148] & !i[1820]) | ( l_42 [8149] &  i[1820]);
assign l_41[6124]    = ( l_42 [8150] & !i[1820]) | ( l_42 [8151] &  i[1820]);
assign l_41[6125]    = ( l_42 [8152] & !i[1820]) | ( l_42 [8153] &  i[1820]);
assign l_41[6126]    = ( l_42 [8154] & !i[1820]) | ( l_42 [8155] &  i[1820]);
assign l_41[6127]    = ( l_42 [8156] & !i[1820]) | ( l_42 [8157] &  i[1820]);
assign l_41[6128]    = ( l_42 [8158] & !i[1820]) | ( l_42 [8159] &  i[1820]);
assign l_41[6129]    = ( l_42 [8160] & !i[1820]) | ( l_42 [8161] &  i[1820]);
assign l_41[6130]    = ( l_42 [8162] & !i[1820]) | ( l_42 [8163] &  i[1820]);
assign l_41[6131]    = ( l_42 [8164] & !i[1820]) | ( l_42 [8165] &  i[1820]);
assign l_41[6132]    = ( l_42 [8166] & !i[1820]) | ( l_42 [8167] &  i[1820]);
assign l_41[6133]    = ( l_42 [8168] & !i[1820]) | ( l_42 [8169] &  i[1820]);
assign l_41[6134]    = ( l_42 [8170] & !i[1820]) | ( l_42 [8171] &  i[1820]);
assign l_41[6135]    = ( l_42 [8172] & !i[1820]) | ( l_42 [8173] &  i[1820]);
assign l_41[6136]    = ( l_42 [8174] & !i[1820]) | ( l_42 [8175] &  i[1820]);
assign l_41[6137]    = ( l_42 [8176] & !i[1820]) | ( l_42 [8177] &  i[1820]);
assign l_41[6138]    = ( l_42 [8178] & !i[1820]) | ( l_42 [8179] &  i[1820]);
assign l_41[6139]    = ( l_42 [8180] & !i[1820]) | ( l_42 [8181] &  i[1820]);
assign l_41[6140]    = ( l_42 [8182] & !i[1820]) | ( l_42 [8183] &  i[1820]);
assign l_41[6141]    = ( l_42 [8184] & !i[1820]) | ( l_42 [8185] &  i[1820]);
assign l_41[6142]    = ( l_42 [8186] & !i[1820]) | ( l_42 [8187] &  i[1820]);
assign l_41[6143]    = ( l_42 [8188] & !i[1820]) | ( l_42 [8189] &  i[1820]);
assign l_41[6144]    = ( l_42 [8190] & !i[1820]) | ( l_42 [8191] &  i[1820]);
assign l_41[6145]    = ( l_42 [8192] & !i[1820]) | ( l_42 [8193] &  i[1820]);
assign l_41[6146]    = ( l_42 [8194] & !i[1820]) | ( l_42 [8195] &  i[1820]);
assign l_41[6147]    = ( l_42 [8196] & !i[1820]) | ( l_42 [8197] &  i[1820]);
assign l_41[6148]    = ( l_42 [8198] & !i[1820]) | ( l_42 [8199] &  i[1820]);
assign l_41[6149]    = ( l_42 [8200] & !i[1820]) | ( l_42 [8201] &  i[1820]);
assign l_41[6150]    = ( l_42 [8202] & !i[1820]) | ( l_42 [8203] &  i[1820]);
assign l_41[6151]    = ( l_42 [8204] & !i[1820]) | ( l_42 [8205] &  i[1820]);
assign l_41[6152]    = ( l_42 [8206] & !i[1820]) | ( l_42 [8207] &  i[1820]);
assign l_41[6153]    = ( l_42 [8208] & !i[1820]) | ( l_42 [8209] &  i[1820]);
assign l_41[6154]    = ( l_42 [8210] & !i[1820]) | ( l_42 [8211] &  i[1820]);
assign l_41[6155]    = ( l_42 [8212] & !i[1820]) | ( l_42 [8213] &  i[1820]);
assign l_41[6156]    = ( l_42 [8214] & !i[1820]) | ( l_42 [8215] &  i[1820]);
assign l_41[6157]    = ( l_42 [8216] & !i[1820]) | ( l_42 [8217] &  i[1820]);
assign l_41[6158]    = ( l_42 [8218] & !i[1820]) | ( l_42 [8219] &  i[1820]);
assign l_41[6159]    = ( l_42 [8220] & !i[1820]) | ( l_42 [8221] &  i[1820]);
assign l_41[6160]    = ( l_42 [8222] & !i[1820]) | ( l_42 [8223] &  i[1820]);
assign l_41[6161]    = ( l_42 [8224] & !i[1820]) | ( l_42 [8225] &  i[1820]);
assign l_41[6162]    = ( l_42 [8226] & !i[1820]) | ( l_42 [8227] &  i[1820]);
assign l_41[6163]    = ( l_42 [8228] & !i[1820]) | ( l_42 [8229] &  i[1820]);
assign l_41[6164]    = ( l_42 [8230] & !i[1820]) | ( l_42 [8231] &  i[1820]);
assign l_41[6165]    = ( l_42 [8232] & !i[1820]) | ( l_42 [8233] &  i[1820]);
assign l_41[6166]    = ( l_42 [8234] & !i[1820]) | ( l_42 [8235] &  i[1820]);
assign l_41[6167]    = ( l_42 [8236] & !i[1820]) | ( l_42 [8237] &  i[1820]);
assign l_41[6168]    = ( l_42 [8238] & !i[1820]) | ( l_42 [8239] &  i[1820]);
assign l_41[6169]    = ( l_42 [8240] & !i[1820]) | ( l_42 [8241] &  i[1820]);
assign l_41[6170]    = ( l_42 [8242] & !i[1820]) | ( l_42 [8243] &  i[1820]);
assign l_41[6171]    = ( l_42 [8244] & !i[1820]) | ( l_42 [8245] &  i[1820]);
assign l_41[6172]    = ( l_42 [8246] & !i[1820]) | ( l_42 [8247] &  i[1820]);
assign l_41[6173]    = ( l_42 [8248] & !i[1820]) | ( l_42 [8249] &  i[1820]);
assign l_41[6174]    = ( l_42 [8250] & !i[1820]) | ( l_42 [8251] &  i[1820]);
assign l_41[6175]    = ( l_42 [8252] & !i[1820]) | ( l_42 [8253] &  i[1820]);
assign l_41[6176]    = ( l_42 [8254] & !i[1820]) | ( l_42 [8255] &  i[1820]);
assign l_41[6177]    = ( l_42 [8256] & !i[1820]) | ( l_42 [8257] &  i[1820]);
assign l_42[0]    = ( l_43 [0] & !i[1703]);
assign l_42[1]    = ( l_43 [1] & !i[1703]) | ( l_43 [2] &  i[1703]);
assign l_42[2]    = ( l_43 [3] & !i[1703]) | ( l_43 [4] &  i[1703]);
assign l_42[3]    = ( l_43 [5] & !i[1703]) | ( l_43 [6] &  i[1703]);
assign l_42[4]    = ( l_43 [7] & !i[1703]) | ( l_43 [8] &  i[1703]);
assign l_42[5]    = ( l_43 [9] & !i[1703]) | ( l_43 [10] &  i[1703]);
assign l_42[6]    = ( l_43 [11] & !i[1703]) | ( l_43 [12] &  i[1703]);
assign l_42[7]    = ( l_43 [13] & !i[1703]) | ( l_43 [14] &  i[1703]);
assign l_42[8]    = ( l_43 [15] & !i[1703]) | ( l_43 [16] &  i[1703]);
assign l_42[9]    = ( l_43 [17] & !i[1703]) | ( l_43 [18] &  i[1703]);
assign l_42[10]    = ( l_43 [19] & !i[1703]) | ( l_43 [20] &  i[1703]);
assign l_42[11]    = ( l_43 [21] & !i[1703]) | ( l_43 [22] &  i[1703]);
assign l_42[12]    = ( l_43 [23] & !i[1703]) | ( l_43 [24] &  i[1703]);
assign l_42[13]    = ( l_43 [25] & !i[1703]) | ( l_43 [26] &  i[1703]);
assign l_42[14]    = ( l_43 [27] & !i[1703]) | ( l_43 [28] &  i[1703]);
assign l_42[15]    = ( l_43 [29] & !i[1703]) | ( l_43 [30] &  i[1703]);
assign l_42[16]    = ( l_43 [31] & !i[1703]) | ( l_43 [32] &  i[1703]);
assign l_42[17]    = ( l_43 [33] & !i[1703]) | ( l_43 [34] &  i[1703]);
assign l_42[18]    = ( l_43 [35] & !i[1703]) | ( l_43 [36] &  i[1703]);
assign l_42[19]    = ( l_43 [37] & !i[1703]) | ( l_43 [38] &  i[1703]);
assign l_42[20]    = ( l_43 [39] & !i[1703]) | ( l_43 [40] &  i[1703]);
assign l_42[21]    = ( l_43 [41] & !i[1703]) | ( l_43 [42] &  i[1703]);
assign l_42[22]    = ( l_43 [43] & !i[1703]) | ( l_43 [44] &  i[1703]);
assign l_42[23]    = ( l_43 [45] & !i[1703]) | ( l_43 [46] &  i[1703]);
assign l_42[24]    = ( l_43 [47] & !i[1703]) | ( l_43 [48] &  i[1703]);
assign l_42[25]    = ( l_43 [49] & !i[1703]) | ( l_43 [50] &  i[1703]);
assign l_42[26]    = ( l_43 [51] & !i[1703]) | ( l_43 [52] &  i[1703]);
assign l_42[27]    = ( l_43 [53] & !i[1703]) | ( l_43 [54] &  i[1703]);
assign l_42[28]    = ( l_43 [55] & !i[1703]) | ( l_43 [56] &  i[1703]);
assign l_42[29]    = ( l_43 [57] & !i[1703]) | ( l_43 [58] &  i[1703]);
assign l_42[30]    = ( l_43 [59] & !i[1703]) | ( l_43 [60] &  i[1703]);
assign l_42[31]    = ( l_43 [61] & !i[1703]) | ( l_43 [62] &  i[1703]);
assign l_42[32]    = ( l_43 [63] & !i[1703]) | ( l_43 [64] &  i[1703]);
assign l_42[33]    = ( l_43 [65] & !i[1703]) | ( l_43 [66] &  i[1703]);
assign l_42[34]    = ( l_43 [67] & !i[1703]) | ( l_43 [68] &  i[1703]);
assign l_42[35]    = ( l_43 [69] & !i[1703]) | ( l_43 [70] &  i[1703]);
assign l_42[36]    = ( l_43 [71] & !i[1703]) | ( l_43 [72] &  i[1703]);
assign l_42[37]    = ( l_43 [73]);
assign l_42[38]    = ( l_43 [74] & !i[1703]) | ( l_43 [75] &  i[1703]);
assign l_42[39]    = ( l_43 [76] & !i[1703]) | ( l_43 [77] &  i[1703]);
assign l_42[40]    = ( l_43 [78] & !i[1703]) | ( l_43 [79] &  i[1703]);
assign l_42[41]    = ( l_43 [80] & !i[1703]) | ( l_43 [81] &  i[1703]);
assign l_42[42]    = ( l_43 [82] & !i[1703]) | ( l_43 [83] &  i[1703]);
assign l_42[43]    = ( l_43 [84] & !i[1703]) | ( l_43 [85] &  i[1703]);
assign l_42[44]    = ( l_43 [86] & !i[1703]) | ( l_43 [87] &  i[1703]);
assign l_42[45]    = ( l_43 [88] & !i[1703]) | ( l_43 [89] &  i[1703]);
assign l_42[46]    = ( l_43 [90] & !i[1703]) | ( l_43 [91] &  i[1703]);
assign l_42[47]    = ( l_43 [92] & !i[1703]) | ( l_43 [93] &  i[1703]);
assign l_42[48]    = ( l_43 [94] & !i[1703]) | ( l_43 [95] &  i[1703]);
assign l_42[49]    = ( l_43 [96] & !i[1703]) | ( l_43 [97] &  i[1703]);
assign l_42[50]    = ( l_43 [98] & !i[1703]) | ( l_43 [99] &  i[1703]);
assign l_42[51]    = ( l_43 [100] & !i[1703]) | ( l_43 [101] &  i[1703]);
assign l_42[52]    = ( l_43 [102] & !i[1703]) | ( l_43 [103] &  i[1703]);
assign l_42[53]    = ( l_43 [104] & !i[1703]) | ( l_43 [105] &  i[1703]);
assign l_42[54]    = ( l_43 [106] & !i[1703]) | ( l_43 [107] &  i[1703]);
assign l_42[55]    = ( l_43 [108] & !i[1703]) | ( l_43 [109] &  i[1703]);
assign l_42[56]    = ( l_43 [110] & !i[1703]) | ( l_43 [111] &  i[1703]);
assign l_42[57]    = ( l_43 [112] & !i[1703]) | ( l_43 [113] &  i[1703]);
assign l_42[58]    = ( l_43 [114] & !i[1703]) | ( l_43 [115] &  i[1703]);
assign l_42[59]    = ( l_43 [116] & !i[1703]) | ( l_43 [117] &  i[1703]);
assign l_42[60]    = ( l_43 [118] & !i[1703]) | ( l_43 [119] &  i[1703]);
assign l_42[61]    = ( l_43 [120] & !i[1703]) | ( l_43 [121] &  i[1703]);
assign l_42[62]    = ( l_43 [122] & !i[1703]) | ( l_43 [123] &  i[1703]);
assign l_42[63]    = ( l_43 [124] & !i[1703]) | ( l_43 [125] &  i[1703]);
assign l_42[64]    = ( l_43 [126] & !i[1703]) | ( l_43 [127] &  i[1703]);
assign l_42[65]    = ( l_43 [128] & !i[1703]) | ( l_43 [129] &  i[1703]);
assign l_42[66]    = ( l_43 [130] & !i[1703]);
assign l_42[67]    = ( l_43 [131] & !i[1703]);
assign l_42[68]    = ( l_43 [132] & !i[1703]);
assign l_42[69]    = ( l_43 [133] & !i[1703]);
assign l_42[70]    = ( l_43 [134] & !i[1703]);
assign l_42[71]    = ( l_43 [135] & !i[1703]);
assign l_42[72]    = ( l_43 [136] & !i[1703]);
assign l_42[73]    = ( l_43 [137] & !i[1703]);
assign l_42[74]    = ( l_43 [130] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[75]    = ( l_43 [131] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[76]    = ( l_43 [132] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[77]    = ( l_43 [133] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[78]    = ( l_43 [134] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[79]    = ( l_43 [135] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[80]    = ( l_43 [136] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[81]    = ( l_43 [137] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[82]    = ( l_43 [130] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[83]    = ( l_43 [131] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[84]    = ( l_43 [132] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[85]    = ( l_43 [133] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[86]    = ( l_43 [134] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[87]    = ( l_43 [135] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[88]    = ( l_43 [136] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[89]    = ( l_43 [137] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[90]    = ( l_43 [130] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[91]    = ( l_43 [131] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[92]    = ( l_43 [132] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[93]    = ( l_43 [133] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[94]    = ( l_43 [134] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[95]    = ( l_43 [135] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[96]    = ( l_43 [136] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[97]    = ( l_43 [137] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[98]    = ( l_43 [130] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[99]    = ( l_43 [131] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[100]    = ( l_43 [132] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[101]    = ( l_43 [133] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[102]    = ( l_43 [134] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[103]    = ( l_43 [135] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[104]    = ( l_43 [136] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[105]    = ( l_43 [137] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[106]    = ( l_43 [130] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[107]    = ( l_43 [131] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[108]    = ( l_43 [132] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[109]    = ( l_43 [133] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[110]    = ( l_43 [134] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[111]    = ( l_43 [135] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[112]    = ( l_43 [136] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[113]    = ( l_43 [137] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[114]    = ( l_43 [130] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[115]    = ( l_43 [131] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[116]    = ( l_43 [132] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[117]    = ( l_43 [133] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[118]    = ( l_43 [134] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[119]    = ( l_43 [135] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[120]    = ( l_43 [136] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[121]    = ( l_43 [137] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[122]    = ( l_43 [130] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[123]    = ( l_43 [131] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[124]    = ( l_43 [132] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[125]    = ( l_43 [133] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[126]    = ( l_43 [134] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[127]    = ( l_43 [135] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[128]    = ( l_43 [136] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[129]    = ( l_43 [137] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[130]    = ( l_43 [130] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[131]    = ( l_43 [131] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[132]    = ( l_43 [132] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[133]    = ( l_43 [133] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[134]    = ( l_43 [134] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[135]    = ( l_43 [135] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[136]    = ( l_43 [136] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[137]    = ( l_43 [137] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[138]    = ( l_43 [130] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[139]    = ( l_43 [131] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[140]    = ( l_43 [132] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[141]    = ( l_43 [133] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[142]    = ( l_43 [134] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[143]    = ( l_43 [135] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[144]    = ( l_43 [136] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[145]    = ( l_43 [137] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[146]    = ( l_43 [130] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[147]    = ( l_43 [131] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[148]    = ( l_43 [132] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[149]    = ( l_43 [133] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[150]    = ( l_43 [134] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[151]    = ( l_43 [135] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[152]    = ( l_43 [136] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[153]    = ( l_43 [137] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[154]    = ( l_43 [130] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[155]    = ( l_43 [131] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[156]    = ( l_43 [132] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[157]    = ( l_43 [133] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[158]    = ( l_43 [134] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[159]    = ( l_43 [135] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[160]    = ( l_43 [136] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[161]    = ( l_43 [137] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[162]    = ( l_43 [130] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[163]    = ( l_43 [131] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[164]    = ( l_43 [132] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[165]    = ( l_43 [133] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[166]    = ( l_43 [134] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[167]    = ( l_43 [135] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[168]    = ( l_43 [136] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[169]    = ( l_43 [137] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[170]    = ( l_43 [130] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[171]    = ( l_43 [131] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[172]    = ( l_43 [132] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[173]    = ( l_43 [133] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[174]    = ( l_43 [134] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[175]    = ( l_43 [135] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[176]    = ( l_43 [136] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[177]    = ( l_43 [137] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[178]    = ( l_43 [130] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[179]    = ( l_43 [131] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[180]    = ( l_43 [132] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[181]    = ( l_43 [133] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[182]    = ( l_43 [134] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[183]    = ( l_43 [135] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[184]    = ( l_43 [136] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[185]    = ( l_43 [137] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[186]    = ( l_43 [130] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[187]    = ( l_43 [131] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[188]    = ( l_43 [132] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[189]    = ( l_43 [133] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[190]    = ( l_43 [134] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[191]    = ( l_43 [135] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[192]    = ( l_43 [136] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[193]    = ( l_43 [137] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[194]    = ( l_43 [130] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[195]    = ( l_43 [131] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[196]    = ( l_43 [132] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[197]    = ( l_43 [133] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[198]    = ( l_43 [134] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[199]    = ( l_43 [135] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[200]    = ( l_43 [136] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[201]    = ( l_43 [137] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[202]    = ( l_43 [130] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[203]    = ( l_43 [131] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[204]    = ( l_43 [132] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[205]    = ( l_43 [133] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[206]    = ( l_43 [134] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[207]    = ( l_43 [135] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[208]    = ( l_43 [136] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[209]    = ( l_43 [137] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[210]    = ( l_43 [130] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[211]    = ( l_43 [131] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[212]    = ( l_43 [132] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[213]    = ( l_43 [133] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[214]    = ( l_43 [134] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[215]    = ( l_43 [135] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[216]    = ( l_43 [136] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[217]    = ( l_43 [137] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[218]    = ( l_43 [130] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[219]    = ( l_43 [131] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[220]    = ( l_43 [132] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[221]    = ( l_43 [133] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[222]    = ( l_43 [134] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[223]    = ( l_43 [135] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[224]    = ( l_43 [136] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[225]    = ( l_43 [137] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[226]    = ( l_43 [130] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[227]    = ( l_43 [131] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[228]    = ( l_43 [132] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[229]    = ( l_43 [133] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[230]    = ( l_43 [134] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[231]    = ( l_43 [135] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[232]    = ( l_43 [136] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[233]    = ( l_43 [137] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[234]    = ( l_43 [130] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[235]    = ( l_43 [131] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[236]    = ( l_43 [132] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[237]    = ( l_43 [133] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[238]    = ( l_43 [134] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[239]    = ( l_43 [135] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[240]    = ( l_43 [136] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[241]    = ( l_43 [137] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[242]    = ( l_43 [130] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[243]    = ( l_43 [131] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[244]    = ( l_43 [132] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[245]    = ( l_43 [133] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[246]    = ( l_43 [134] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[247]    = ( l_43 [135] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[248]    = ( l_43 [136] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[249]    = ( l_43 [137] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[250]    = ( l_43 [130] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[251]    = ( l_43 [131] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[252]    = ( l_43 [132] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[253]    = ( l_43 [133] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[254]    = ( l_43 [134] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[255]    = ( l_43 [135] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[256]    = ( l_43 [136] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[257]    = ( l_43 [137] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[258]    = ( l_43 [130] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[259]    = ( l_43 [131] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[260]    = ( l_43 [132] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[261]    = ( l_43 [133] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[262]    = ( l_43 [134] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[263]    = ( l_43 [135] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[264]    = ( l_43 [136] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[265]    = ( l_43 [137] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[266]    = ( l_43 [130] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[267]    = ( l_43 [131] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[268]    = ( l_43 [132] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[269]    = ( l_43 [133] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[270]    = ( l_43 [134] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[271]    = ( l_43 [135] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[272]    = ( l_43 [136] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[273]    = ( l_43 [137] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[274]    = ( l_43 [130] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[275]    = ( l_43 [131] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[276]    = ( l_43 [132] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[277]    = ( l_43 [133] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[278]    = ( l_43 [134] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[279]    = ( l_43 [135] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[280]    = ( l_43 [136] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[281]    = ( l_43 [137] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[282]    = ( l_43 [130] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[283]    = ( l_43 [131] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[284]    = ( l_43 [132] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[285]    = ( l_43 [133] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[286]    = ( l_43 [134] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[287]    = ( l_43 [135] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[288]    = ( l_43 [136] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[289]    = ( l_43 [137] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[290]    = ( l_43 [130] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[291]    = ( l_43 [131] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[292]    = ( l_43 [132] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[293]    = ( l_43 [133] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[294]    = ( l_43 [134] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[295]    = ( l_43 [135] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[296]    = ( l_43 [136] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[297]    = ( l_43 [137] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[298]    = ( l_43 [130] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[299]    = ( l_43 [131] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[300]    = ( l_43 [132] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[301]    = ( l_43 [133] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[302]    = ( l_43 [134] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[303]    = ( l_43 [135] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[304]    = ( l_43 [136] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[305]    = ( l_43 [137] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[306]    = ( l_43 [130] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[307]    = ( l_43 [131] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[308]    = ( l_43 [132] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[309]    = ( l_43 [133] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[310]    = ( l_43 [134] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[311]    = ( l_43 [135] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[312]    = ( l_43 [136] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[313]    = ( l_43 [137] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[314]    = ( l_43 [130] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[315]    = ( l_43 [131] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[316]    = ( l_43 [132] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[317]    = ( l_43 [133] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[318]    = ( l_43 [134] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[319]    = ( l_43 [135] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[320]    = ( l_43 [136] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[321]    = ( l_43 [137] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[322]    = ( l_43 [130] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[323]    = ( l_43 [131] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[324]    = ( l_43 [132] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[325]    = ( l_43 [133] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[326]    = ( l_43 [134] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[327]    = ( l_43 [135] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[328]    = ( l_43 [136] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[329]    = ( l_43 [137] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[330]    = ( l_43 [130] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[331]    = ( l_43 [131] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[332]    = ( l_43 [132] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[333]    = ( l_43 [133] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[334]    = ( l_43 [134] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[335]    = ( l_43 [135] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[336]    = ( l_43 [136] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[337]    = ( l_43 [137] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[338]    = ( l_43 [130] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[339]    = ( l_43 [131] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[340]    = ( l_43 [132] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[341]    = ( l_43 [133] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[342]    = ( l_43 [134] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[343]    = ( l_43 [135] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[344]    = ( l_43 [136] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[345]    = ( l_43 [137] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[346]    = ( l_43 [130] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[347]    = ( l_43 [131] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[348]    = ( l_43 [132] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[349]    = ( l_43 [133] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[350]    = ( l_43 [134] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[351]    = ( l_43 [135] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[352]    = ( l_43 [136] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[353]    = ( l_43 [137] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[354]    = ( l_43 [130] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[355]    = ( l_43 [131] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[356]    = ( l_43 [132] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[357]    = ( l_43 [133] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[358]    = ( l_43 [134] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[359]    = ( l_43 [135] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[360]    = ( l_43 [136] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[361]    = ( l_43 [137] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[362]    = ( l_43 [130] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[363]    = ( l_43 [131] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[364]    = ( l_43 [132] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[365]    = ( l_43 [133] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[366]    = ( l_43 [134] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[367]    = ( l_43 [135] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[368]    = ( l_43 [136] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[369]    = ( l_43 [137] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[370]    = ( l_43 [130] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[371]    = ( l_43 [131] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[372]    = ( l_43 [132] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[373]    = ( l_43 [133] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[374]    = ( l_43 [134] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[375]    = ( l_43 [135] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[376]    = ( l_43 [136] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[377]    = ( l_43 [137] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[378]    = ( l_43 [130] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[379]    = ( l_43 [131] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[380]    = ( l_43 [132] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[381]    = ( l_43 [133] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[382]    = ( l_43 [134] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[383]    = ( l_43 [135] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[384]    = ( l_43 [136] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[385]    = ( l_43 [137] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[386]    = ( l_43 [130] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[387]    = ( l_43 [131] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[388]    = ( l_43 [132] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[389]    = ( l_43 [133] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[390]    = ( l_43 [134] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[391]    = ( l_43 [135] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[392]    = ( l_43 [136] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[393]    = ( l_43 [137] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[394]    = ( l_43 [130] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[395]    = ( l_43 [131] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[396]    = ( l_43 [132] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[397]    = ( l_43 [133] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[398]    = ( l_43 [134] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[399]    = ( l_43 [135] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[400]    = ( l_43 [136] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[401]    = ( l_43 [137] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[402]    = ( l_43 [130] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[403]    = ( l_43 [131] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[404]    = ( l_43 [132] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[405]    = ( l_43 [133] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[406]    = ( l_43 [134] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[407]    = ( l_43 [135] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[408]    = ( l_43 [136] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[409]    = ( l_43 [137] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[410]    = ( l_43 [130] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[411]    = ( l_43 [131] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[412]    = ( l_43 [132] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[413]    = ( l_43 [133] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[414]    = ( l_43 [134] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[415]    = ( l_43 [135] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[416]    = ( l_43 [136] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[417]    = ( l_43 [137] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[418]    = ( l_43 [130] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[419]    = ( l_43 [131] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[420]    = ( l_43 [132] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[421]    = ( l_43 [133] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[422]    = ( l_43 [134] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[423]    = ( l_43 [135] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[424]    = ( l_43 [136] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[425]    = ( l_43 [137] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[426]    = ( l_43 [130] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[427]    = ( l_43 [131] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[428]    = ( l_43 [132] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[429]    = ( l_43 [133] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[430]    = ( l_43 [134] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[431]    = ( l_43 [135] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[432]    = ( l_43 [136] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[433]    = ( l_43 [137] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[434]    = ( l_43 [130] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[435]    = ( l_43 [131] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[436]    = ( l_43 [132] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[437]    = ( l_43 [133] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[438]    = ( l_43 [134] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[439]    = ( l_43 [135] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[440]    = ( l_43 [136] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[441]    = ( l_43 [137] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[442]    = ( l_43 [130] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[443]    = ( l_43 [131] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[444]    = ( l_43 [132] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[445]    = ( l_43 [133] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[446]    = ( l_43 [134] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[447]    = ( l_43 [135] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[448]    = ( l_43 [136] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[449]    = ( l_43 [137] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[450]    = ( l_43 [130] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[451]    = ( l_43 [131] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[452]    = ( l_43 [132] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[453]    = ( l_43 [133] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[454]    = ( l_43 [134] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[455]    = ( l_43 [135] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[456]    = ( l_43 [136] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[457]    = ( l_43 [137] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[458]    = ( l_43 [130] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[459]    = ( l_43 [131] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[460]    = ( l_43 [132] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[461]    = ( l_43 [133] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[462]    = ( l_43 [134] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[463]    = ( l_43 [135] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[464]    = ( l_43 [136] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[465]    = ( l_43 [137] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[466]    = ( l_43 [130] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[467]    = ( l_43 [131] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[468]    = ( l_43 [132] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[469]    = ( l_43 [133] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[470]    = ( l_43 [134] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[471]    = ( l_43 [135] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[472]    = ( l_43 [136] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[473]    = ( l_43 [137] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[474]    = ( l_43 [130] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[475]    = ( l_43 [131] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[476]    = ( l_43 [132] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[477]    = ( l_43 [133] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[478]    = ( l_43 [134] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[479]    = ( l_43 [135] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[480]    = ( l_43 [136] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[481]    = ( l_43 [137] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[482]    = ( l_43 [130] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[483]    = ( l_43 [131] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[484]    = ( l_43 [132] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[485]    = ( l_43 [133] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[486]    = ( l_43 [134] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[487]    = ( l_43 [135] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[488]    = ( l_43 [136] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[489]    = ( l_43 [137] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[490]    = ( l_43 [130] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[491]    = ( l_43 [131] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[492]    = ( l_43 [132] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[493]    = ( l_43 [133] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[494]    = ( l_43 [134] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[495]    = ( l_43 [135] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[496]    = ( l_43 [136] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[497]    = ( l_43 [137] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[498]    = ( l_43 [130] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[499]    = ( l_43 [131] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[500]    = ( l_43 [132] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[501]    = ( l_43 [133] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[502]    = ( l_43 [134] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[503]    = ( l_43 [135] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[504]    = ( l_43 [136] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[505]    = ( l_43 [137] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[506]    = ( l_43 [130] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[507]    = ( l_43 [131] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[508]    = ( l_43 [132] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[509]    = ( l_43 [133] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[510]    = ( l_43 [134] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[511]    = ( l_43 [135] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[512]    = ( l_43 [136] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[513]    = ( l_43 [137] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[514]    = ( l_43 [130] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[515]    = ( l_43 [131] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[516]    = ( l_43 [132] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[517]    = ( l_43 [133] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[518]    = ( l_43 [134] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[519]    = ( l_43 [135] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[520]    = ( l_43 [136] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[521]    = ( l_43 [137] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[522]    = ( l_43 [130] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[523]    = ( l_43 [131] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[524]    = ( l_43 [132] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[525]    = ( l_43 [133] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[526]    = ( l_43 [134] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[527]    = ( l_43 [135] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[528]    = ( l_43 [136] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[529]    = ( l_43 [137] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[530]    = ( l_43 [130] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[531]    = ( l_43 [131] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[532]    = ( l_43 [132] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[533]    = ( l_43 [133] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[534]    = ( l_43 [134] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[535]    = ( l_43 [135] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[536]    = ( l_43 [136] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[537]    = ( l_43 [137] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[538]    = ( l_43 [130] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[539]    = ( l_43 [131] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[540]    = ( l_43 [132] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[541]    = ( l_43 [133] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[542]    = ( l_43 [134] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[543]    = ( l_43 [135] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[544]    = ( l_43 [136] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[545]    = ( l_43 [137] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[546]    = ( l_43 [130] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[547]    = ( l_43 [131] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[548]    = ( l_43 [132] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[549]    = ( l_43 [133] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[550]    = ( l_43 [134] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[551]    = ( l_43 [135] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[552]    = ( l_43 [136] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[553]    = ( l_43 [137] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[554]    = ( l_43 [130] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[555]    = ( l_43 [131] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[556]    = ( l_43 [132] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[557]    = ( l_43 [133] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[558]    = ( l_43 [134] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[559]    = ( l_43 [135] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[560]    = ( l_43 [136] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[561]    = ( l_43 [137] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[562]    = ( l_43 [130] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[563]    = ( l_43 [131] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[564]    = ( l_43 [132] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[565]    = ( l_43 [133] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[566]    = ( l_43 [134] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[567]    = ( l_43 [135] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[568]    = ( l_43 [136] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[569]    = ( l_43 [137] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[570]    = ( l_43 [130] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[571]    = ( l_43 [131] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[572]    = ( l_43 [132] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[573]    = ( l_43 [133] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[574]    = ( l_43 [134] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[575]    = ( l_43 [135] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[576]    = ( l_43 [136] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[577]    = ( l_43 [137] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[578]    = ( l_43 [130] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[579]    = ( l_43 [131] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[580]    = ( l_43 [132] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[581]    = ( l_43 [133] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[582]    = ( l_43 [134] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[583]    = ( l_43 [135] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[584]    = ( l_43 [136] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[585]    = ( l_43 [137] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[586]    = ( l_43 [130] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[587]    = ( l_43 [131] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[588]    = ( l_43 [132] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[589]    = ( l_43 [133] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[590]    = ( l_43 [134] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[591]    = ( l_43 [135] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[592]    = ( l_43 [136] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[593]    = ( l_43 [137] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[594]    = ( l_43 [130] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[595]    = ( l_43 [131] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[596]    = ( l_43 [132] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[597]    = ( l_43 [133] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[598]    = ( l_43 [134] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[599]    = ( l_43 [135] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[600]    = ( l_43 [136] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[601]    = ( l_43 [137] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[602]    = ( l_43 [130] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[603]    = ( l_43 [131] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[604]    = ( l_43 [132] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[605]    = ( l_43 [133] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[606]    = ( l_43 [134] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[607]    = ( l_43 [135] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[608]    = ( l_43 [136] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[609]    = ( l_43 [137] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[610]    = ( l_43 [130] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[611]    = ( l_43 [131] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[612]    = ( l_43 [132] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[613]    = ( l_43 [133] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[614]    = ( l_43 [134] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[615]    = ( l_43 [135] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[616]    = ( l_43 [136] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[617]    = ( l_43 [137] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[618]    = ( l_43 [130] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[619]    = ( l_43 [131] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[620]    = ( l_43 [132] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[621]    = ( l_43 [133] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[622]    = ( l_43 [134] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[623]    = ( l_43 [135] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[624]    = ( l_43 [136] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[625]    = ( l_43 [137] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[626]    = ( l_43 [130] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[627]    = ( l_43 [131] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[628]    = ( l_43 [132] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[629]    = ( l_43 [133] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[630]    = ( l_43 [134] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[631]    = ( l_43 [135] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[632]    = ( l_43 [136] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[633]    = ( l_43 [137] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[634]    = ( l_43 [130] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[635]    = ( l_43 [131] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[636]    = ( l_43 [132] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[637]    = ( l_43 [133] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[638]    = ( l_43 [134] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[639]    = ( l_43 [135] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[640]    = ( l_43 [136] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[641]    = ( l_43 [137] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[642]    = ( l_43 [130] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[643]    = ( l_43 [131] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[644]    = ( l_43 [132] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[645]    = ( l_43 [133] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[646]    = ( l_43 [134] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[647]    = ( l_43 [135] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[648]    = ( l_43 [136] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[649]    = ( l_43 [137] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[650]    = ( l_43 [130] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[651]    = ( l_43 [131] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[652]    = ( l_43 [132] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[653]    = ( l_43 [133] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[654]    = ( l_43 [134] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[655]    = ( l_43 [135] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[656]    = ( l_43 [136] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[657]    = ( l_43 [137] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[658]    = ( l_43 [130] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[659]    = ( l_43 [131] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[660]    = ( l_43 [132] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[661]    = ( l_43 [133] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[662]    = ( l_43 [134] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[663]    = ( l_43 [135] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[664]    = ( l_43 [136] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[665]    = ( l_43 [137] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[666]    = ( l_43 [130] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[667]    = ( l_43 [131] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[668]    = ( l_43 [132] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[669]    = ( l_43 [133] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[670]    = ( l_43 [134] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[671]    = ( l_43 [135] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[672]    = ( l_43 [136] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[673]    = ( l_43 [137] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[674]    = ( l_43 [130] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[675]    = ( l_43 [131] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[676]    = ( l_43 [132] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[677]    = ( l_43 [133] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[678]    = ( l_43 [134] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[679]    = ( l_43 [135] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[680]    = ( l_43 [136] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[681]    = ( l_43 [137] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[682]    = ( l_43 [130] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[683]    = ( l_43 [131] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[684]    = ( l_43 [132] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[685]    = ( l_43 [133] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[686]    = ( l_43 [134] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[687]    = ( l_43 [135] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[688]    = ( l_43 [136] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[689]    = ( l_43 [137] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[690]    = ( l_43 [130] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[691]    = ( l_43 [131] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[692]    = ( l_43 [132] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[693]    = ( l_43 [133] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[694]    = ( l_43 [134] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[695]    = ( l_43 [135] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[696]    = ( l_43 [136] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[697]    = ( l_43 [137] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[698]    = ( l_43 [130] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[699]    = ( l_43 [131] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[700]    = ( l_43 [132] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[701]    = ( l_43 [133] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[702]    = ( l_43 [134] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[703]    = ( l_43 [135] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[704]    = ( l_43 [136] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[705]    = ( l_43 [137] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[706]    = ( l_43 [130] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[707]    = ( l_43 [131] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[708]    = ( l_43 [132] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[709]    = ( l_43 [133] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[710]    = ( l_43 [134] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[711]    = ( l_43 [135] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[712]    = ( l_43 [136] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[713]    = ( l_43 [137] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[714]    = ( l_43 [130] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[715]    = ( l_43 [131] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[716]    = ( l_43 [132] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[717]    = ( l_43 [133] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[718]    = ( l_43 [134] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[719]    = ( l_43 [135] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[720]    = ( l_43 [136] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[721]    = ( l_43 [137] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[722]    = ( l_43 [130] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[723]    = ( l_43 [131] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[724]    = ( l_43 [132] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[725]    = ( l_43 [133] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[726]    = ( l_43 [134] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[727]    = ( l_43 [135] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[728]    = ( l_43 [136] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[729]    = ( l_43 [137] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[730]    = ( l_43 [130] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[731]    = ( l_43 [131] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[732]    = ( l_43 [132] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[733]    = ( l_43 [133] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[734]    = ( l_43 [134] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[735]    = ( l_43 [135] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[736]    = ( l_43 [136] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[737]    = ( l_43 [137] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[738]    = ( l_43 [130] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[739]    = ( l_43 [131] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[740]    = ( l_43 [132] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[741]    = ( l_43 [133] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[742]    = ( l_43 [134] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[743]    = ( l_43 [135] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[744]    = ( l_43 [136] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[745]    = ( l_43 [137] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[746]    = ( l_43 [130] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[747]    = ( l_43 [131] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[748]    = ( l_43 [132] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[749]    = ( l_43 [133] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[750]    = ( l_43 [134] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[751]    = ( l_43 [135] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[752]    = ( l_43 [136] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[753]    = ( l_43 [137] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[754]    = ( l_43 [130] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[755]    = ( l_43 [131] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[756]    = ( l_43 [132] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[757]    = ( l_43 [133] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[758]    = ( l_43 [134] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[759]    = ( l_43 [135] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[760]    = ( l_43 [136] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[761]    = ( l_43 [137] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[762]    = ( l_43 [130] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[763]    = ( l_43 [131] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[764]    = ( l_43 [132] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[765]    = ( l_43 [133] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[766]    = ( l_43 [134] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[767]    = ( l_43 [135] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[768]    = ( l_43 [136] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[769]    = ( l_43 [137] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[770]    = ( l_43 [130] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[771]    = ( l_43 [131] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[772]    = ( l_43 [132] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[773]    = ( l_43 [133] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[774]    = ( l_43 [134] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[775]    = ( l_43 [135] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[776]    = ( l_43 [136] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[777]    = ( l_43 [137] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[778]    = ( l_43 [130] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[779]    = ( l_43 [131] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[780]    = ( l_43 [132] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[781]    = ( l_43 [133] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[782]    = ( l_43 [134] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[783]    = ( l_43 [135] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[784]    = ( l_43 [136] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[785]    = ( l_43 [137] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[786]    = ( l_43 [130] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[787]    = ( l_43 [131] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[788]    = ( l_43 [132] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[789]    = ( l_43 [133] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[790]    = ( l_43 [134] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[791]    = ( l_43 [135] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[792]    = ( l_43 [136] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[793]    = ( l_43 [137] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[794]    = ( l_43 [130] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[795]    = ( l_43 [131] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[796]    = ( l_43 [132] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[797]    = ( l_43 [133] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[798]    = ( l_43 [134] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[799]    = ( l_43 [135] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[800]    = ( l_43 [136] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[801]    = ( l_43 [137] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[802]    = ( l_43 [130] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[803]    = ( l_43 [131] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[804]    = ( l_43 [132] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[805]    = ( l_43 [133] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[806]    = ( l_43 [134] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[807]    = ( l_43 [135] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[808]    = ( l_43 [136] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[809]    = ( l_43 [137] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[810]    = ( l_43 [130] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[811]    = ( l_43 [131] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[812]    = ( l_43 [132] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[813]    = ( l_43 [133] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[814]    = ( l_43 [134] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[815]    = ( l_43 [135] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[816]    = ( l_43 [136] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[817]    = ( l_43 [137] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[818]    = ( l_43 [130] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[819]    = ( l_43 [131] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[820]    = ( l_43 [132] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[821]    = ( l_43 [133] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[822]    = ( l_43 [134] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[823]    = ( l_43 [135] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[824]    = ( l_43 [136] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[825]    = ( l_43 [137] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[826]    = ( l_43 [130] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[827]    = ( l_43 [131] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[828]    = ( l_43 [132] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[829]    = ( l_43 [133] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[830]    = ( l_43 [134] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[831]    = ( l_43 [135] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[832]    = ( l_43 [136] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[833]    = ( l_43 [137] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[834]    = ( l_43 [130] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[835]    = ( l_43 [131] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[836]    = ( l_43 [132] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[837]    = ( l_43 [133] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[838]    = ( l_43 [134] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[839]    = ( l_43 [135] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[840]    = ( l_43 [136] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[841]    = ( l_43 [137] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[842]    = ( l_43 [130] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[843]    = ( l_43 [131] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[844]    = ( l_43 [132] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[845]    = ( l_43 [133] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[846]    = ( l_43 [134] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[847]    = ( l_43 [135] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[848]    = ( l_43 [136] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[849]    = ( l_43 [137] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[850]    = ( l_43 [130] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[851]    = ( l_43 [131] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[852]    = ( l_43 [132] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[853]    = ( l_43 [133] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[854]    = ( l_43 [134] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[855]    = ( l_43 [135] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[856]    = ( l_43 [136] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[857]    = ( l_43 [137] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[858]    = ( l_43 [130] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[859]    = ( l_43 [131] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[860]    = ( l_43 [132] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[861]    = ( l_43 [133] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[862]    = ( l_43 [134] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[863]    = ( l_43 [135] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[864]    = ( l_43 [136] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[865]    = ( l_43 [137] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[866]    = ( l_43 [130] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[867]    = ( l_43 [131] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[868]    = ( l_43 [132] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[869]    = ( l_43 [133] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[870]    = ( l_43 [134] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[871]    = ( l_43 [135] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[872]    = ( l_43 [136] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[873]    = ( l_43 [137] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[874]    = ( l_43 [130] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[875]    = ( l_43 [131] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[876]    = ( l_43 [132] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[877]    = ( l_43 [133] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[878]    = ( l_43 [134] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[879]    = ( l_43 [135] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[880]    = ( l_43 [136] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[881]    = ( l_43 [137] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[882]    = ( l_43 [130] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[883]    = ( l_43 [131] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[884]    = ( l_43 [132] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[885]    = ( l_43 [133] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[886]    = ( l_43 [134] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[887]    = ( l_43 [135] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[888]    = ( l_43 [136] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[889]    = ( l_43 [137] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[890]    = ( l_43 [130] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[891]    = ( l_43 [131] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[892]    = ( l_43 [132] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[893]    = ( l_43 [133] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[894]    = ( l_43 [134] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[895]    = ( l_43 [135] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[896]    = ( l_43 [136] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[897]    = ( l_43 [137] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[898]    = ( l_43 [130] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[899]    = ( l_43 [131] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[900]    = ( l_43 [132] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[901]    = ( l_43 [133] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[902]    = ( l_43 [134] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[903]    = ( l_43 [135] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[904]    = ( l_43 [136] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[905]    = ( l_43 [137] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[906]    = ( l_43 [130] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[907]    = ( l_43 [131] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[908]    = ( l_43 [132] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[909]    = ( l_43 [133] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[910]    = ( l_43 [134] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[911]    = ( l_43 [135] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[912]    = ( l_43 [136] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[913]    = ( l_43 [137] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[914]    = ( l_43 [130] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[915]    = ( l_43 [131] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[916]    = ( l_43 [132] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[917]    = ( l_43 [133] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[918]    = ( l_43 [134] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[919]    = ( l_43 [135] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[920]    = ( l_43 [136] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[921]    = ( l_43 [137] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[922]    = ( l_43 [130] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[923]    = ( l_43 [131] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[924]    = ( l_43 [132] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[925]    = ( l_43 [133] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[926]    = ( l_43 [134] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[927]    = ( l_43 [135] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[928]    = ( l_43 [136] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[929]    = ( l_43 [137] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[930]    = ( l_43 [130] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[931]    = ( l_43 [131] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[932]    = ( l_43 [132] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[933]    = ( l_43 [133] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[934]    = ( l_43 [134] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[935]    = ( l_43 [135] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[936]    = ( l_43 [136] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[937]    = ( l_43 [137] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[938]    = ( l_43 [130] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[939]    = ( l_43 [131] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[940]    = ( l_43 [132] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[941]    = ( l_43 [133] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[942]    = ( l_43 [134] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[943]    = ( l_43 [135] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[944]    = ( l_43 [136] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[945]    = ( l_43 [137] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[946]    = ( l_43 [130] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[947]    = ( l_43 [131] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[948]    = ( l_43 [132] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[949]    = ( l_43 [133] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[950]    = ( l_43 [134] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[951]    = ( l_43 [135] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[952]    = ( l_43 [136] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[953]    = ( l_43 [137] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[954]    = ( l_43 [130] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[955]    = ( l_43 [131] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[956]    = ( l_43 [132] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[957]    = ( l_43 [133] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[958]    = ( l_43 [134] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[959]    = ( l_43 [135] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[960]    = ( l_43 [136] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[961]    = ( l_43 [137] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[962]    = ( l_43 [130] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[963]    = ( l_43 [131] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[964]    = ( l_43 [132] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[965]    = ( l_43 [133] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[966]    = ( l_43 [134] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[967]    = ( l_43 [135] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[968]    = ( l_43 [136] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[969]    = ( l_43 [137] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[970]    = ( l_43 [130] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[971]    = ( l_43 [131] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[972]    = ( l_43 [132] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[973]    = ( l_43 [133] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[974]    = ( l_43 [134] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[975]    = ( l_43 [135] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[976]    = ( l_43 [136] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[977]    = ( l_43 [137] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[978]    = ( l_43 [130] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[979]    = ( l_43 [131] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[980]    = ( l_43 [132] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[981]    = ( l_43 [133] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[982]    = ( l_43 [134] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[983]    = ( l_43 [135] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[984]    = ( l_43 [136] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[985]    = ( l_43 [137] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[986]    = ( l_43 [130] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[987]    = ( l_43 [131] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[988]    = ( l_43 [132] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[989]    = ( l_43 [133] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[990]    = ( l_43 [134] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[991]    = ( l_43 [135] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[992]    = ( l_43 [136] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[993]    = ( l_43 [137] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[994]    = ( l_43 [130] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[995]    = ( l_43 [131] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[996]    = ( l_43 [132] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[997]    = ( l_43 [133] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[998]    = ( l_43 [134] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[999]    = ( l_43 [135] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[1000]    = ( l_43 [136] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[1001]    = ( l_43 [137] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[1002]    = ( l_43 [130] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1003]    = ( l_43 [131] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1004]    = ( l_43 [132] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1005]    = ( l_43 [133] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1006]    = ( l_43 [134] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1007]    = ( l_43 [135] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1008]    = ( l_43 [136] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1009]    = ( l_43 [137] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[1010]    = ( l_43 [130] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1011]    = ( l_43 [131] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1012]    = ( l_43 [132] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1013]    = ( l_43 [133] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1014]    = ( l_43 [134] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1015]    = ( l_43 [135] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1016]    = ( l_43 [136] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1017]    = ( l_43 [137] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[1018]    = ( l_43 [130] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1019]    = ( l_43 [131] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1020]    = ( l_43 [132] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1021]    = ( l_43 [133] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1022]    = ( l_43 [134] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1023]    = ( l_43 [135] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1024]    = ( l_43 [136] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1025]    = ( l_43 [137] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[1026]    = ( l_43 [130] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1027]    = ( l_43 [131] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1028]    = ( l_43 [132] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1029]    = ( l_43 [133] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1030]    = ( l_43 [134] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1031]    = ( l_43 [135] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1032]    = ( l_43 [136] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1033]    = ( l_43 [137] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[1034]    = ( l_43 [130] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1035]    = ( l_43 [131] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1036]    = ( l_43 [132] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1037]    = ( l_43 [133] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1038]    = ( l_43 [134] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1039]    = ( l_43 [135] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1040]    = ( l_43 [136] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1041]    = ( l_43 [137] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[1042]    = ( l_43 [130] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1043]    = ( l_43 [131] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1044]    = ( l_43 [132] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1045]    = ( l_43 [133] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1046]    = ( l_43 [134] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1047]    = ( l_43 [135] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1048]    = ( l_43 [136] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1049]    = ( l_43 [137] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[1050]    = ( l_43 [130] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1051]    = ( l_43 [131] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1052]    = ( l_43 [132] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1053]    = ( l_43 [133] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1054]    = ( l_43 [134] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1055]    = ( l_43 [135] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1056]    = ( l_43 [136] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1057]    = ( l_43 [137] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[1058]    = ( l_43 [130] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1059]    = ( l_43 [131] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1060]    = ( l_43 [132] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1061]    = ( l_43 [133] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1062]    = ( l_43 [134] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1063]    = ( l_43 [135] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1064]    = ( l_43 [136] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1065]    = ( l_43 [137] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[1066]    = ( l_43 [130] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1067]    = ( l_43 [131] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1068]    = ( l_43 [132] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1069]    = ( l_43 [133] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1070]    = ( l_43 [134] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1071]    = ( l_43 [135] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1072]    = ( l_43 [136] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1073]    = ( l_43 [137] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[1074]    = ( l_43 [130] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1075]    = ( l_43 [131] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1076]    = ( l_43 [132] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1077]    = ( l_43 [133] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1078]    = ( l_43 [134] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1079]    = ( l_43 [135] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1080]    = ( l_43 [136] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1081]    = ( l_43 [137] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[1082]    = ( l_43 [130] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1083]    = ( l_43 [131] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1084]    = ( l_43 [132] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1085]    = ( l_43 [133] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1086]    = ( l_43 [134] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1087]    = ( l_43 [135] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1088]    = ( l_43 [136] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1089]    = ( l_43 [137] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[1090]    = ( l_43 [130] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1091]    = ( l_43 [131] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1092]    = ( l_43 [132] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1093]    = ( l_43 [133] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1094]    = ( l_43 [134] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1095]    = ( l_43 [135] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1096]    = ( l_43 [136] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1097]    = ( l_43 [137] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[1098]    = ( l_43 [130] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1099]    = ( l_43 [131] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1100]    = ( l_43 [132] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1101]    = ( l_43 [133] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1102]    = ( l_43 [134] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1103]    = ( l_43 [135] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1104]    = ( l_43 [136] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1105]    = ( l_43 [137] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[1106]    = ( l_43 [130] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1107]    = ( l_43 [131] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1108]    = ( l_43 [132] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1109]    = ( l_43 [133] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1110]    = ( l_43 [134] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1111]    = ( l_43 [135] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1112]    = ( l_43 [136] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1113]    = ( l_43 [137] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[1114]    = ( l_43 [130] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1115]    = ( l_43 [131] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1116]    = ( l_43 [132] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1117]    = ( l_43 [133] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1118]    = ( l_43 [134] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1119]    = ( l_43 [135] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1120]    = ( l_43 [136] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1121]    = ( l_43 [137] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[1122]    = ( l_43 [130] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1123]    = ( l_43 [131] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1124]    = ( l_43 [132] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1125]    = ( l_43 [133] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1126]    = ( l_43 [134] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1127]    = ( l_43 [135] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1128]    = ( l_43 [136] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1129]    = ( l_43 [137] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[1130]    = ( l_43 [130] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1131]    = ( l_43 [131] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1132]    = ( l_43 [132] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1133]    = ( l_43 [133] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1134]    = ( l_43 [134] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1135]    = ( l_43 [135] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1136]    = ( l_43 [136] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1137]    = ( l_43 [137] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[1138]    = ( l_43 [130] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1139]    = ( l_43 [131] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1140]    = ( l_43 [132] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1141]    = ( l_43 [133] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1142]    = ( l_43 [134] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1143]    = ( l_43 [135] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1144]    = ( l_43 [136] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1145]    = ( l_43 [137] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[1146]    = ( l_43 [130] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1147]    = ( l_43 [131] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1148]    = ( l_43 [132] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1149]    = ( l_43 [133] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1150]    = ( l_43 [134] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1151]    = ( l_43 [135] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1152]    = ( l_43 [136] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1153]    = ( l_43 [137] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[1154]    = ( l_43 [130] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1155]    = ( l_43 [131] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1156]    = ( l_43 [132] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1157]    = ( l_43 [133] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1158]    = ( l_43 [134] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1159]    = ( l_43 [135] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1160]    = ( l_43 [136] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1161]    = ( l_43 [137] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[1162]    = ( l_43 [130] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1163]    = ( l_43 [131] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1164]    = ( l_43 [132] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1165]    = ( l_43 [133] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1166]    = ( l_43 [134] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1167]    = ( l_43 [135] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1168]    = ( l_43 [136] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1169]    = ( l_43 [137] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[1170]    = ( l_43 [130] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1171]    = ( l_43 [131] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1172]    = ( l_43 [132] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1173]    = ( l_43 [133] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1174]    = ( l_43 [134] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1175]    = ( l_43 [135] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1176]    = ( l_43 [136] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1177]    = ( l_43 [137] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[1178]    = ( l_43 [130] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1179]    = ( l_43 [131] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1180]    = ( l_43 [132] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1181]    = ( l_43 [133] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1182]    = ( l_43 [134] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1183]    = ( l_43 [135] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1184]    = ( l_43 [136] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1185]    = ( l_43 [137] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[1186]    = ( l_43 [130] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1187]    = ( l_43 [131] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1188]    = ( l_43 [132] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1189]    = ( l_43 [133] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1190]    = ( l_43 [134] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1191]    = ( l_43 [135] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1192]    = ( l_43 [136] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1193]    = ( l_43 [137] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[1194]    = ( l_43 [130] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1195]    = ( l_43 [131] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1196]    = ( l_43 [132] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1197]    = ( l_43 [133] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1198]    = ( l_43 [134] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1199]    = ( l_43 [135] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1200]    = ( l_43 [136] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1201]    = ( l_43 [137] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[1202]    = ( l_43 [130] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1203]    = ( l_43 [131] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1204]    = ( l_43 [132] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1205]    = ( l_43 [133] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1206]    = ( l_43 [134] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1207]    = ( l_43 [135] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1208]    = ( l_43 [136] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1209]    = ( l_43 [137] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[1210]    = ( l_43 [130] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1211]    = ( l_43 [131] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1212]    = ( l_43 [132] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1213]    = ( l_43 [133] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1214]    = ( l_43 [134] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1215]    = ( l_43 [135] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1216]    = ( l_43 [136] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1217]    = ( l_43 [137] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[1218]    = ( l_43 [130] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1219]    = ( l_43 [131] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1220]    = ( l_43 [132] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1221]    = ( l_43 [133] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1222]    = ( l_43 [134] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1223]    = ( l_43 [135] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1224]    = ( l_43 [136] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1225]    = ( l_43 [137] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[1226]    = ( l_43 [130] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1227]    = ( l_43 [131] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1228]    = ( l_43 [132] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1229]    = ( l_43 [133] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1230]    = ( l_43 [134] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1231]    = ( l_43 [135] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1232]    = ( l_43 [136] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1233]    = ( l_43 [137] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[1234]    = ( l_43 [130] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1235]    = ( l_43 [131] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1236]    = ( l_43 [132] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1237]    = ( l_43 [133] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1238]    = ( l_43 [134] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1239]    = ( l_43 [135] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1240]    = ( l_43 [136] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1241]    = ( l_43 [137] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[1242]    = ( l_43 [130] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1243]    = ( l_43 [131] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1244]    = ( l_43 [132] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1245]    = ( l_43 [133] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1246]    = ( l_43 [134] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1247]    = ( l_43 [135] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1248]    = ( l_43 [136] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1249]    = ( l_43 [137] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[1250]    = ( l_43 [130] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1251]    = ( l_43 [131] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1252]    = ( l_43 [132] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1253]    = ( l_43 [133] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1254]    = ( l_43 [134] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1255]    = ( l_43 [135] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1256]    = ( l_43 [136] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1257]    = ( l_43 [137] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[1258]    = ( l_43 [130] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1259]    = ( l_43 [131] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1260]    = ( l_43 [132] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1261]    = ( l_43 [133] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1262]    = ( l_43 [134] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1263]    = ( l_43 [135] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1264]    = ( l_43 [136] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1265]    = ( l_43 [137] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[1266]    = ( l_43 [130] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1267]    = ( l_43 [131] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1268]    = ( l_43 [132] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1269]    = ( l_43 [133] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1270]    = ( l_43 [134] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1271]    = ( l_43 [135] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1272]    = ( l_43 [136] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1273]    = ( l_43 [137] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[1274]    = ( l_43 [130] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1275]    = ( l_43 [131] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1276]    = ( l_43 [132] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1277]    = ( l_43 [133] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1278]    = ( l_43 [134] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1279]    = ( l_43 [135] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1280]    = ( l_43 [136] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1281]    = ( l_43 [137] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[1282]    = ( l_43 [130] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1283]    = ( l_43 [131] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1284]    = ( l_43 [132] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1285]    = ( l_43 [133] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1286]    = ( l_43 [134] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1287]    = ( l_43 [135] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1288]    = ( l_43 [136] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1289]    = ( l_43 [137] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[1290]    = ( l_43 [130] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1291]    = ( l_43 [131] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1292]    = ( l_43 [132] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1293]    = ( l_43 [133] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1294]    = ( l_43 [134] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1295]    = ( l_43 [135] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1296]    = ( l_43 [136] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1297]    = ( l_43 [137] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[1298]    = ( l_43 [130] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1299]    = ( l_43 [131] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1300]    = ( l_43 [132] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1301]    = ( l_43 [133] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1302]    = ( l_43 [134] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1303]    = ( l_43 [135] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1304]    = ( l_43 [136] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1305]    = ( l_43 [137] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[1306]    = ( l_43 [130] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1307]    = ( l_43 [131] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1308]    = ( l_43 [132] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1309]    = ( l_43 [133] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1310]    = ( l_43 [134] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1311]    = ( l_43 [135] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1312]    = ( l_43 [136] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1313]    = ( l_43 [137] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[1314]    = ( l_43 [130] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1315]    = ( l_43 [131] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1316]    = ( l_43 [132] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1317]    = ( l_43 [133] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1318]    = ( l_43 [134] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1319]    = ( l_43 [135] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1320]    = ( l_43 [136] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1321]    = ( l_43 [137] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[1322]    = ( l_43 [130] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1323]    = ( l_43 [131] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1324]    = ( l_43 [132] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1325]    = ( l_43 [133] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1326]    = ( l_43 [134] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1327]    = ( l_43 [135] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1328]    = ( l_43 [136] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1329]    = ( l_43 [137] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[1330]    = ( l_43 [130] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1331]    = ( l_43 [131] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1332]    = ( l_43 [132] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1333]    = ( l_43 [133] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1334]    = ( l_43 [134] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1335]    = ( l_43 [135] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1336]    = ( l_43 [136] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1337]    = ( l_43 [137] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[1338]    = ( l_43 [130] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1339]    = ( l_43 [131] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1340]    = ( l_43 [132] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1341]    = ( l_43 [133] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1342]    = ( l_43 [134] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1343]    = ( l_43 [135] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1344]    = ( l_43 [136] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1345]    = ( l_43 [137] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[1346]    = ( l_43 [130] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1347]    = ( l_43 [131] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1348]    = ( l_43 [132] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1349]    = ( l_43 [133] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1350]    = ( l_43 [134] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1351]    = ( l_43 [135] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1352]    = ( l_43 [136] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1353]    = ( l_43 [137] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[1354]    = ( l_43 [130] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1355]    = ( l_43 [131] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1356]    = ( l_43 [132] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1357]    = ( l_43 [133] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1358]    = ( l_43 [134] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1359]    = ( l_43 [135] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1360]    = ( l_43 [136] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1361]    = ( l_43 [137] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[1362]    = ( l_43 [130] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1363]    = ( l_43 [131] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1364]    = ( l_43 [132] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1365]    = ( l_43 [133] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1366]    = ( l_43 [134] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1367]    = ( l_43 [135] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1368]    = ( l_43 [136] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1369]    = ( l_43 [137] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[1370]    = ( l_43 [130] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1371]    = ( l_43 [131] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1372]    = ( l_43 [132] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1373]    = ( l_43 [133] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1374]    = ( l_43 [134] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1375]    = ( l_43 [135] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1376]    = ( l_43 [136] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1377]    = ( l_43 [137] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[1378]    = ( l_43 [130] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1379]    = ( l_43 [131] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1380]    = ( l_43 [132] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1381]    = ( l_43 [133] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1382]    = ( l_43 [134] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1383]    = ( l_43 [135] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1384]    = ( l_43 [136] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1385]    = ( l_43 [137] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[1386]    = ( l_43 [130] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1387]    = ( l_43 [131] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1388]    = ( l_43 [132] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1389]    = ( l_43 [133] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1390]    = ( l_43 [134] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1391]    = ( l_43 [135] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1392]    = ( l_43 [136] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1393]    = ( l_43 [137] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[1394]    = ( l_43 [130] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1395]    = ( l_43 [131] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1396]    = ( l_43 [132] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1397]    = ( l_43 [133] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1398]    = ( l_43 [134] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1399]    = ( l_43 [135] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1400]    = ( l_43 [136] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1401]    = ( l_43 [137] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[1402]    = ( l_43 [130] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1403]    = ( l_43 [131] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1404]    = ( l_43 [132] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1405]    = ( l_43 [133] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1406]    = ( l_43 [134] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1407]    = ( l_43 [135] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1408]    = ( l_43 [136] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1409]    = ( l_43 [137] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[1410]    = ( l_43 [130] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1411]    = ( l_43 [131] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1412]    = ( l_43 [132] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1413]    = ( l_43 [133] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1414]    = ( l_43 [134] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1415]    = ( l_43 [135] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1416]    = ( l_43 [136] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1417]    = ( l_43 [137] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[1418]    = ( l_43 [130] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1419]    = ( l_43 [131] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1420]    = ( l_43 [132] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1421]    = ( l_43 [133] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1422]    = ( l_43 [134] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1423]    = ( l_43 [135] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1424]    = ( l_43 [136] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1425]    = ( l_43 [137] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[1426]    = ( l_43 [130] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1427]    = ( l_43 [131] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1428]    = ( l_43 [132] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1429]    = ( l_43 [133] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1430]    = ( l_43 [134] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1431]    = ( l_43 [135] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1432]    = ( l_43 [136] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1433]    = ( l_43 [137] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[1434]    = ( l_43 [130] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1435]    = ( l_43 [131] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1436]    = ( l_43 [132] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1437]    = ( l_43 [133] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1438]    = ( l_43 [134] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1439]    = ( l_43 [135] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1440]    = ( l_43 [136] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1441]    = ( l_43 [137] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[1442]    = ( l_43 [130] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1443]    = ( l_43 [131] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1444]    = ( l_43 [132] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1445]    = ( l_43 [133] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1446]    = ( l_43 [134] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1447]    = ( l_43 [135] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1448]    = ( l_43 [136] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1449]    = ( l_43 [137] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[1450]    = ( l_43 [130] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1451]    = ( l_43 [131] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1452]    = ( l_43 [132] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1453]    = ( l_43 [133] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1454]    = ( l_43 [134] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1455]    = ( l_43 [135] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1456]    = ( l_43 [136] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1457]    = ( l_43 [137] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[1458]    = ( l_43 [130] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1459]    = ( l_43 [131] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1460]    = ( l_43 [132] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1461]    = ( l_43 [133] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1462]    = ( l_43 [134] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1463]    = ( l_43 [135] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1464]    = ( l_43 [136] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1465]    = ( l_43 [137] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[1466]    = ( l_43 [130] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1467]    = ( l_43 [131] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1468]    = ( l_43 [132] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1469]    = ( l_43 [133] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1470]    = ( l_43 [134] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1471]    = ( l_43 [135] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1472]    = ( l_43 [136] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1473]    = ( l_43 [137] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[1474]    = ( l_43 [130] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1475]    = ( l_43 [131] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1476]    = ( l_43 [132] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1477]    = ( l_43 [133] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1478]    = ( l_43 [134] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1479]    = ( l_43 [135] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1480]    = ( l_43 [136] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1481]    = ( l_43 [137] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[1482]    = ( l_43 [130] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1483]    = ( l_43 [131] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1484]    = ( l_43 [132] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1485]    = ( l_43 [133] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1486]    = ( l_43 [134] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1487]    = ( l_43 [135] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1488]    = ( l_43 [136] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1489]    = ( l_43 [137] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[1490]    = ( l_43 [130] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1491]    = ( l_43 [131] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1492]    = ( l_43 [132] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1493]    = ( l_43 [133] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1494]    = ( l_43 [134] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1495]    = ( l_43 [135] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1496]    = ( l_43 [136] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1497]    = ( l_43 [137] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[1498]    = ( l_43 [130] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1499]    = ( l_43 [131] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1500]    = ( l_43 [132] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1501]    = ( l_43 [133] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1502]    = ( l_43 [134] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1503]    = ( l_43 [135] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1504]    = ( l_43 [136] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1505]    = ( l_43 [137] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[1506]    = ( l_43 [130] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1507]    = ( l_43 [131] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1508]    = ( l_43 [132] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1509]    = ( l_43 [133] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1510]    = ( l_43 [134] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1511]    = ( l_43 [135] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1512]    = ( l_43 [136] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1513]    = ( l_43 [137] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[1514]    = ( l_43 [130] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1515]    = ( l_43 [131] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1516]    = ( l_43 [132] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1517]    = ( l_43 [133] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1518]    = ( l_43 [134] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1519]    = ( l_43 [135] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1520]    = ( l_43 [136] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1521]    = ( l_43 [137] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[1522]    = ( l_43 [130] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1523]    = ( l_43 [131] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1524]    = ( l_43 [132] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1525]    = ( l_43 [133] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1526]    = ( l_43 [134] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1527]    = ( l_43 [135] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1528]    = ( l_43 [136] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1529]    = ( l_43 [137] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[1530]    = ( l_43 [130] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1531]    = ( l_43 [131] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1532]    = ( l_43 [132] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1533]    = ( l_43 [133] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1534]    = ( l_43 [134] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1535]    = ( l_43 [135] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1536]    = ( l_43 [136] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1537]    = ( l_43 [137] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[1538]    = ( l_43 [130] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1539]    = ( l_43 [131] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1540]    = ( l_43 [132] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1541]    = ( l_43 [133] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1542]    = ( l_43 [134] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1543]    = ( l_43 [135] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1544]    = ( l_43 [136] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1545]    = ( l_43 [137] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[1546]    = ( l_43 [130] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1547]    = ( l_43 [131] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1548]    = ( l_43 [132] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1549]    = ( l_43 [133] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1550]    = ( l_43 [134] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1551]    = ( l_43 [135] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1552]    = ( l_43 [136] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1553]    = ( l_43 [137] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[1554]    = ( l_43 [130] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1555]    = ( l_43 [131] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1556]    = ( l_43 [132] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1557]    = ( l_43 [133] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1558]    = ( l_43 [134] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1559]    = ( l_43 [135] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1560]    = ( l_43 [136] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1561]    = ( l_43 [137] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[1562]    = ( l_43 [130] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1563]    = ( l_43 [131] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1564]    = ( l_43 [132] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1565]    = ( l_43 [133] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1566]    = ( l_43 [134] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1567]    = ( l_43 [135] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1568]    = ( l_43 [136] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1569]    = ( l_43 [137] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[1570]    = ( l_43 [130] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1571]    = ( l_43 [131] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1572]    = ( l_43 [132] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1573]    = ( l_43 [133] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1574]    = ( l_43 [134] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1575]    = ( l_43 [135] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1576]    = ( l_43 [136] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1577]    = ( l_43 [137] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[1578]    = ( l_43 [130] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1579]    = ( l_43 [131] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1580]    = ( l_43 [132] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1581]    = ( l_43 [133] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1582]    = ( l_43 [134] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1583]    = ( l_43 [135] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1584]    = ( l_43 [136] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1585]    = ( l_43 [137] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[1586]    = ( l_43 [130] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1587]    = ( l_43 [131] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1588]    = ( l_43 [132] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1589]    = ( l_43 [133] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1590]    = ( l_43 [134] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1591]    = ( l_43 [135] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1592]    = ( l_43 [136] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1593]    = ( l_43 [137] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[1594]    = ( l_43 [130] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1595]    = ( l_43 [131] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1596]    = ( l_43 [132] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1597]    = ( l_43 [133] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1598]    = ( l_43 [134] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1599]    = ( l_43 [135] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1600]    = ( l_43 [136] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1601]    = ( l_43 [137] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[1602]    = ( l_43 [130] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1603]    = ( l_43 [131] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1604]    = ( l_43 [132] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1605]    = ( l_43 [133] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1606]    = ( l_43 [134] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1607]    = ( l_43 [135] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1608]    = ( l_43 [136] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1609]    = ( l_43 [137] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[1610]    = ( l_43 [130] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1611]    = ( l_43 [131] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1612]    = ( l_43 [132] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1613]    = ( l_43 [133] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1614]    = ( l_43 [134] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1615]    = ( l_43 [135] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1616]    = ( l_43 [136] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1617]    = ( l_43 [137] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[1618]    = ( l_43 [130] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1619]    = ( l_43 [131] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1620]    = ( l_43 [132] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1621]    = ( l_43 [133] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1622]    = ( l_43 [134] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1623]    = ( l_43 [135] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1624]    = ( l_43 [136] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1625]    = ( l_43 [137] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[1626]    = ( l_43 [130] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1627]    = ( l_43 [131] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1628]    = ( l_43 [132] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1629]    = ( l_43 [133] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1630]    = ( l_43 [134] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1631]    = ( l_43 [135] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1632]    = ( l_43 [136] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1633]    = ( l_43 [137] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[1634]    = ( l_43 [130] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1635]    = ( l_43 [131] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1636]    = ( l_43 [132] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1637]    = ( l_43 [133] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1638]    = ( l_43 [134] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1639]    = ( l_43 [135] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1640]    = ( l_43 [136] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1641]    = ( l_43 [137] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[1642]    = ( l_43 [130] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1643]    = ( l_43 [131] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1644]    = ( l_43 [132] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1645]    = ( l_43 [133] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1646]    = ( l_43 [134] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1647]    = ( l_43 [135] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1648]    = ( l_43 [136] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1649]    = ( l_43 [137] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[1650]    = ( l_43 [130] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1651]    = ( l_43 [131] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1652]    = ( l_43 [132] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1653]    = ( l_43 [133] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1654]    = ( l_43 [134] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1655]    = ( l_43 [135] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1656]    = ( l_43 [136] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1657]    = ( l_43 [137] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[1658]    = ( l_43 [130] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1659]    = ( l_43 [131] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1660]    = ( l_43 [132] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1661]    = ( l_43 [133] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1662]    = ( l_43 [134] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1663]    = ( l_43 [135] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1664]    = ( l_43 [136] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1665]    = ( l_43 [137] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[1666]    = ( l_43 [130] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1667]    = ( l_43 [131] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1668]    = ( l_43 [132] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1669]    = ( l_43 [133] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1670]    = ( l_43 [134] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1671]    = ( l_43 [135] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1672]    = ( l_43 [136] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1673]    = ( l_43 [137] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[1674]    = ( l_43 [130] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1675]    = ( l_43 [131] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1676]    = ( l_43 [132] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1677]    = ( l_43 [133] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1678]    = ( l_43 [134] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1679]    = ( l_43 [135] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1680]    = ( l_43 [136] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1681]    = ( l_43 [137] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[1682]    = ( l_43 [130] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1683]    = ( l_43 [131] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1684]    = ( l_43 [132] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1685]    = ( l_43 [133] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1686]    = ( l_43 [134] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1687]    = ( l_43 [135] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1688]    = ( l_43 [136] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1689]    = ( l_43 [137] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[1690]    = ( l_43 [130] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1691]    = ( l_43 [131] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1692]    = ( l_43 [132] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1693]    = ( l_43 [133] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1694]    = ( l_43 [134] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1695]    = ( l_43 [135] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1696]    = ( l_43 [136] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1697]    = ( l_43 [137] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[1698]    = ( l_43 [130] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1699]    = ( l_43 [131] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1700]    = ( l_43 [132] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1701]    = ( l_43 [133] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1702]    = ( l_43 [134] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1703]    = ( l_43 [135] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1704]    = ( l_43 [136] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1705]    = ( l_43 [137] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[1706]    = ( l_43 [130] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1707]    = ( l_43 [131] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1708]    = ( l_43 [132] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1709]    = ( l_43 [133] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1710]    = ( l_43 [134] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1711]    = ( l_43 [135] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1712]    = ( l_43 [136] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1713]    = ( l_43 [137] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[1714]    = ( l_43 [130] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1715]    = ( l_43 [131] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1716]    = ( l_43 [132] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1717]    = ( l_43 [133] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1718]    = ( l_43 [134] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1719]    = ( l_43 [135] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1720]    = ( l_43 [136] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1721]    = ( l_43 [137] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[1722]    = ( l_43 [130] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1723]    = ( l_43 [131] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1724]    = ( l_43 [132] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1725]    = ( l_43 [133] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1726]    = ( l_43 [134] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1727]    = ( l_43 [135] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1728]    = ( l_43 [136] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1729]    = ( l_43 [137] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[1730]    = ( l_43 [130] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1731]    = ( l_43 [131] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1732]    = ( l_43 [132] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1733]    = ( l_43 [133] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1734]    = ( l_43 [134] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1735]    = ( l_43 [135] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1736]    = ( l_43 [136] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1737]    = ( l_43 [137] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[1738]    = ( l_43 [130] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1739]    = ( l_43 [131] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1740]    = ( l_43 [132] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1741]    = ( l_43 [133] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1742]    = ( l_43 [134] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1743]    = ( l_43 [135] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1744]    = ( l_43 [136] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1745]    = ( l_43 [137] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[1746]    = ( l_43 [130] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1747]    = ( l_43 [131] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1748]    = ( l_43 [132] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1749]    = ( l_43 [133] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1750]    = ( l_43 [134] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1751]    = ( l_43 [135] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1752]    = ( l_43 [136] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1753]    = ( l_43 [137] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[1754]    = ( l_43 [130] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1755]    = ( l_43 [131] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1756]    = ( l_43 [132] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1757]    = ( l_43 [133] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1758]    = ( l_43 [134] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1759]    = ( l_43 [135] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1760]    = ( l_43 [136] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1761]    = ( l_43 [137] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[1762]    = ( l_43 [130] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1763]    = ( l_43 [131] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1764]    = ( l_43 [132] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1765]    = ( l_43 [133] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1766]    = ( l_43 [134] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1767]    = ( l_43 [135] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1768]    = ( l_43 [136] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1769]    = ( l_43 [137] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[1770]    = ( l_43 [130] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1771]    = ( l_43 [131] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1772]    = ( l_43 [132] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1773]    = ( l_43 [133] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1774]    = ( l_43 [134] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1775]    = ( l_43 [135] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1776]    = ( l_43 [136] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1777]    = ( l_43 [137] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[1778]    = ( l_43 [130] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1779]    = ( l_43 [131] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1780]    = ( l_43 [132] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1781]    = ( l_43 [133] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1782]    = ( l_43 [134] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1783]    = ( l_43 [135] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1784]    = ( l_43 [136] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1785]    = ( l_43 [137] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[1786]    = ( l_43 [130] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1787]    = ( l_43 [131] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1788]    = ( l_43 [132] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1789]    = ( l_43 [133] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1790]    = ( l_43 [134] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1791]    = ( l_43 [135] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1792]    = ( l_43 [136] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1793]    = ( l_43 [137] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[1794]    = ( l_43 [130] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1795]    = ( l_43 [131] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1796]    = ( l_43 [132] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1797]    = ( l_43 [133] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1798]    = ( l_43 [134] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1799]    = ( l_43 [135] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1800]    = ( l_43 [136] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1801]    = ( l_43 [137] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[1802]    = ( l_43 [130] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1803]    = ( l_43 [131] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1804]    = ( l_43 [132] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1805]    = ( l_43 [133] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1806]    = ( l_43 [134] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1807]    = ( l_43 [135] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1808]    = ( l_43 [136] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1809]    = ( l_43 [137] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[1810]    = ( l_43 [130] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1811]    = ( l_43 [131] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1812]    = ( l_43 [132] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1813]    = ( l_43 [133] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1814]    = ( l_43 [134] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1815]    = ( l_43 [135] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1816]    = ( l_43 [136] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1817]    = ( l_43 [137] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[1818]    = ( l_43 [130] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1819]    = ( l_43 [131] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1820]    = ( l_43 [132] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1821]    = ( l_43 [133] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1822]    = ( l_43 [134] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1823]    = ( l_43 [135] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1824]    = ( l_43 [136] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1825]    = ( l_43 [137] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[1826]    = ( l_43 [130] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1827]    = ( l_43 [131] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1828]    = ( l_43 [132] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1829]    = ( l_43 [133] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1830]    = ( l_43 [134] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1831]    = ( l_43 [135] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1832]    = ( l_43 [136] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1833]    = ( l_43 [137] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[1834]    = ( l_43 [130] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1835]    = ( l_43 [131] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1836]    = ( l_43 [132] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1837]    = ( l_43 [133] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1838]    = ( l_43 [134] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1839]    = ( l_43 [135] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1840]    = ( l_43 [136] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1841]    = ( l_43 [137] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[1842]    = ( l_43 [130] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1843]    = ( l_43 [131] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1844]    = ( l_43 [132] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1845]    = ( l_43 [133] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1846]    = ( l_43 [134] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1847]    = ( l_43 [135] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1848]    = ( l_43 [136] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1849]    = ( l_43 [137] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[1850]    = ( l_43 [130] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1851]    = ( l_43 [131] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1852]    = ( l_43 [132] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1853]    = ( l_43 [133] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1854]    = ( l_43 [134] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1855]    = ( l_43 [135] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1856]    = ( l_43 [136] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1857]    = ( l_43 [137] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[1858]    = ( l_43 [130] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1859]    = ( l_43 [131] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1860]    = ( l_43 [132] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1861]    = ( l_43 [133] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1862]    = ( l_43 [134] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1863]    = ( l_43 [135] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1864]    = ( l_43 [136] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1865]    = ( l_43 [137] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[1866]    = ( l_43 [130] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1867]    = ( l_43 [131] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1868]    = ( l_43 [132] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1869]    = ( l_43 [133] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1870]    = ( l_43 [134] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1871]    = ( l_43 [135] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1872]    = ( l_43 [136] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1873]    = ( l_43 [137] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[1874]    = ( l_43 [130] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1875]    = ( l_43 [131] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1876]    = ( l_43 [132] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1877]    = ( l_43 [133] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1878]    = ( l_43 [134] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1879]    = ( l_43 [135] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1880]    = ( l_43 [136] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1881]    = ( l_43 [137] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[1882]    = ( l_43 [130] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1883]    = ( l_43 [131] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1884]    = ( l_43 [132] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1885]    = ( l_43 [133] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1886]    = ( l_43 [134] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1887]    = ( l_43 [135] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1888]    = ( l_43 [136] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1889]    = ( l_43 [137] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[1890]    = ( l_43 [130] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1891]    = ( l_43 [131] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1892]    = ( l_43 [132] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1893]    = ( l_43 [133] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1894]    = ( l_43 [134] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1895]    = ( l_43 [135] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1896]    = ( l_43 [136] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1897]    = ( l_43 [137] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[1898]    = ( l_43 [130] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1899]    = ( l_43 [131] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1900]    = ( l_43 [132] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1901]    = ( l_43 [133] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1902]    = ( l_43 [134] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1903]    = ( l_43 [135] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1904]    = ( l_43 [136] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1905]    = ( l_43 [137] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[1906]    = ( l_43 [130] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1907]    = ( l_43 [131] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1908]    = ( l_43 [132] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1909]    = ( l_43 [133] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1910]    = ( l_43 [134] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1911]    = ( l_43 [135] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1912]    = ( l_43 [136] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1913]    = ( l_43 [137] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[1914]    = ( l_43 [130] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1915]    = ( l_43 [131] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1916]    = ( l_43 [132] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1917]    = ( l_43 [133] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1918]    = ( l_43 [134] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1919]    = ( l_43 [135] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1920]    = ( l_43 [136] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1921]    = ( l_43 [137] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[1922]    = ( l_43 [130] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1923]    = ( l_43 [131] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1924]    = ( l_43 [132] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1925]    = ( l_43 [133] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1926]    = ( l_43 [134] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1927]    = ( l_43 [135] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1928]    = ( l_43 [136] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1929]    = ( l_43 [137] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[1930]    = ( l_43 [130] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1931]    = ( l_43 [131] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1932]    = ( l_43 [132] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1933]    = ( l_43 [133] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1934]    = ( l_43 [134] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1935]    = ( l_43 [135] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1936]    = ( l_43 [136] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1937]    = ( l_43 [137] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[1938]    = ( l_43 [130] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1939]    = ( l_43 [131] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1940]    = ( l_43 [132] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1941]    = ( l_43 [133] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1942]    = ( l_43 [134] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1943]    = ( l_43 [135] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1944]    = ( l_43 [136] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1945]    = ( l_43 [137] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[1946]    = ( l_43 [130] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1947]    = ( l_43 [131] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1948]    = ( l_43 [132] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1949]    = ( l_43 [133] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1950]    = ( l_43 [134] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1951]    = ( l_43 [135] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1952]    = ( l_43 [136] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1953]    = ( l_43 [137] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[1954]    = ( l_43 [130] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1955]    = ( l_43 [131] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1956]    = ( l_43 [132] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1957]    = ( l_43 [133] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1958]    = ( l_43 [134] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1959]    = ( l_43 [135] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1960]    = ( l_43 [136] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1961]    = ( l_43 [137] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[1962]    = ( l_43 [130] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1963]    = ( l_43 [131] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1964]    = ( l_43 [132] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1965]    = ( l_43 [133] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1966]    = ( l_43 [134] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1967]    = ( l_43 [135] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1968]    = ( l_43 [136] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1969]    = ( l_43 [137] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[1970]    = ( l_43 [130] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1971]    = ( l_43 [131] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1972]    = ( l_43 [132] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1973]    = ( l_43 [133] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1974]    = ( l_43 [134] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1975]    = ( l_43 [135] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1976]    = ( l_43 [136] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1977]    = ( l_43 [137] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[1978]    = ( l_43 [130] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1979]    = ( l_43 [131] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1980]    = ( l_43 [132] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1981]    = ( l_43 [133] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1982]    = ( l_43 [134] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1983]    = ( l_43 [135] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1984]    = ( l_43 [136] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1985]    = ( l_43 [137] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[1986]    = ( l_43 [130] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1987]    = ( l_43 [131] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1988]    = ( l_43 [132] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1989]    = ( l_43 [133] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1990]    = ( l_43 [134] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1991]    = ( l_43 [135] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1992]    = ( l_43 [136] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1993]    = ( l_43 [137] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[1994]    = ( l_43 [130] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[1995]    = ( l_43 [131] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[1996]    = ( l_43 [132] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[1997]    = ( l_43 [133] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[1998]    = ( l_43 [134] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[1999]    = ( l_43 [135] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[2000]    = ( l_43 [136] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[2001]    = ( l_43 [137] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[2002]    = ( l_43 [130] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2003]    = ( l_43 [131] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2004]    = ( l_43 [132] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2005]    = ( l_43 [133] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2006]    = ( l_43 [134] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2007]    = ( l_43 [135] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2008]    = ( l_43 [136] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2009]    = ( l_43 [137] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[2010]    = ( l_43 [130] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2011]    = ( l_43 [131] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2012]    = ( l_43 [132] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2013]    = ( l_43 [133] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2014]    = ( l_43 [134] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2015]    = ( l_43 [135] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2016]    = ( l_43 [136] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2017]    = ( l_43 [137] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[2018]    = ( l_43 [130] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2019]    = ( l_43 [131] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2020]    = ( l_43 [132] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2021]    = ( l_43 [133] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2022]    = ( l_43 [134] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2023]    = ( l_43 [135] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2024]    = ( l_43 [136] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2025]    = ( l_43 [137] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[2026]    = ( l_43 [130] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2027]    = ( l_43 [131] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2028]    = ( l_43 [132] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2029]    = ( l_43 [133] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2030]    = ( l_43 [134] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2031]    = ( l_43 [135] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2032]    = ( l_43 [136] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2033]    = ( l_43 [137] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[2034]    = ( l_43 [130] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2035]    = ( l_43 [131] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2036]    = ( l_43 [132] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2037]    = ( l_43 [133] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2038]    = ( l_43 [134] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2039]    = ( l_43 [135] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2040]    = ( l_43 [136] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2041]    = ( l_43 [137] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[2042]    = ( l_43 [130] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2043]    = ( l_43 [131] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2044]    = ( l_43 [132] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2045]    = ( l_43 [133] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2046]    = ( l_43 [134] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2047]    = ( l_43 [135] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2048]    = ( l_43 [136] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2049]    = ( l_43 [137] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[2050]    = ( l_43 [130] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2051]    = ( l_43 [131] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2052]    = ( l_43 [132] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2053]    = ( l_43 [133] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2054]    = ( l_43 [134] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2055]    = ( l_43 [135] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2056]    = ( l_43 [136] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2057]    = ( l_43 [137] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[2058]    = ( l_43 [130] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2059]    = ( l_43 [131] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2060]    = ( l_43 [132] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2061]    = ( l_43 [133] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2062]    = ( l_43 [134] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2063]    = ( l_43 [135] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2064]    = ( l_43 [136] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2065]    = ( l_43 [137] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[2066]    = ( l_43 [130] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2067]    = ( l_43 [131] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2068]    = ( l_43 [132] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2069]    = ( l_43 [133] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2070]    = ( l_43 [134] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2071]    = ( l_43 [135] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2072]    = ( l_43 [136] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2073]    = ( l_43 [137] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[2074]    = ( l_43 [130] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2075]    = ( l_43 [131] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2076]    = ( l_43 [132] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2077]    = ( l_43 [133] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2078]    = ( l_43 [134] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2079]    = ( l_43 [135] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2080]    = ( l_43 [136] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2081]    = ( l_43 [137] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[2082]    = ( l_43 [130] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2083]    = ( l_43 [131] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2084]    = ( l_43 [132] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2085]    = ( l_43 [133] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2086]    = ( l_43 [134] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2087]    = ( l_43 [135] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2088]    = ( l_43 [136] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2089]    = ( l_43 [137] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[2090]    = ( l_43 [130] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2091]    = ( l_43 [131] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2092]    = ( l_43 [132] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2093]    = ( l_43 [133] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2094]    = ( l_43 [134] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2095]    = ( l_43 [135] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2096]    = ( l_43 [136] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2097]    = ( l_43 [137] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[2098]    = ( l_43 [130] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2099]    = ( l_43 [131] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2100]    = ( l_43 [132] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2101]    = ( l_43 [133] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2102]    = ( l_43 [134] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2103]    = ( l_43 [135] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2104]    = ( l_43 [136] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2105]    = ( l_43 [137] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[2106]    = ( l_43 [130] & !i[1703]) | (      i[1703]);
assign l_42[2107]    = ( l_43 [131] & !i[1703]) | (      i[1703]);
assign l_42[2108]    = ( l_43 [132] & !i[1703]) | (      i[1703]);
assign l_42[2109]    = ( l_43 [133] & !i[1703]) | (      i[1703]);
assign l_42[2110]    = ( l_43 [134] & !i[1703]) | (      i[1703]);
assign l_42[2111]    = ( l_43 [135] & !i[1703]) | (      i[1703]);
assign l_42[2112]    = ( l_43 [136] & !i[1703]) | (      i[1703]);
assign l_42[2113]    = ( l_43 [137] & !i[1703]) | (      i[1703]);
assign l_42[2114]    = ( l_43 [391] & !i[1703]);
assign l_42[2115]    = ( l_43 [392] & !i[1703]);
assign l_42[2116]    = ( l_43 [393] & !i[1703]);
assign l_42[2117]    = ( l_43 [394] & !i[1703]);
assign l_42[2118]    = ( l_43 [395] & !i[1703]);
assign l_42[2119]    = ( l_43 [396] & !i[1703]);
assign l_42[2120]    = ( l_43 [397] & !i[1703]);
assign l_42[2121]    = ( l_43 [398] & !i[1703]);
assign l_42[2122]    = ( l_43 [391] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2123]    = ( l_43 [392] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2124]    = ( l_43 [393] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2125]    = ( l_43 [394] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2126]    = ( l_43 [395] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2127]    = ( l_43 [396] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2128]    = ( l_43 [397] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2129]    = ( l_43 [398] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[2130]    = ( l_43 [391] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2131]    = ( l_43 [392] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2132]    = ( l_43 [393] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2133]    = ( l_43 [394] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2134]    = ( l_43 [395] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2135]    = ( l_43 [396] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2136]    = ( l_43 [397] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2137]    = ( l_43 [398] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[2138]    = ( l_43 [391] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2139]    = ( l_43 [392] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2140]    = ( l_43 [393] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2141]    = ( l_43 [394] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2142]    = ( l_43 [395] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2143]    = ( l_43 [396] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2144]    = ( l_43 [397] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2145]    = ( l_43 [398] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[2146]    = ( l_43 [391] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2147]    = ( l_43 [392] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2148]    = ( l_43 [393] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2149]    = ( l_43 [394] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2150]    = ( l_43 [395] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2151]    = ( l_43 [396] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2152]    = ( l_43 [397] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2153]    = ( l_43 [398] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[2154]    = ( l_43 [391] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2155]    = ( l_43 [392] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2156]    = ( l_43 [393] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2157]    = ( l_43 [394] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2158]    = ( l_43 [395] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2159]    = ( l_43 [396] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2160]    = ( l_43 [397] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2161]    = ( l_43 [398] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[2162]    = ( l_43 [391] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2163]    = ( l_43 [392] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2164]    = ( l_43 [393] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2165]    = ( l_43 [394] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2166]    = ( l_43 [395] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2167]    = ( l_43 [396] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2168]    = ( l_43 [397] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2169]    = ( l_43 [398] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[2170]    = ( l_43 [391] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2171]    = ( l_43 [392] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2172]    = ( l_43 [393] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2173]    = ( l_43 [394] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2174]    = ( l_43 [395] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2175]    = ( l_43 [396] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2176]    = ( l_43 [397] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2177]    = ( l_43 [398] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[2178]    = ( l_43 [391] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2179]    = ( l_43 [392] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2180]    = ( l_43 [393] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2181]    = ( l_43 [394] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2182]    = ( l_43 [395] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2183]    = ( l_43 [396] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2184]    = ( l_43 [397] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2185]    = ( l_43 [398] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[2186]    = ( l_43 [391] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2187]    = ( l_43 [392] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2188]    = ( l_43 [393] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2189]    = ( l_43 [394] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2190]    = ( l_43 [395] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2191]    = ( l_43 [396] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2192]    = ( l_43 [397] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2193]    = ( l_43 [398] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[2194]    = ( l_43 [391] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2195]    = ( l_43 [392] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2196]    = ( l_43 [393] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2197]    = ( l_43 [394] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2198]    = ( l_43 [395] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2199]    = ( l_43 [396] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2200]    = ( l_43 [397] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2201]    = ( l_43 [398] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[2202]    = ( l_43 [391] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2203]    = ( l_43 [392] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2204]    = ( l_43 [393] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2205]    = ( l_43 [394] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2206]    = ( l_43 [395] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2207]    = ( l_43 [396] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2208]    = ( l_43 [397] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2209]    = ( l_43 [398] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[2210]    = ( l_43 [391] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2211]    = ( l_43 [392] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2212]    = ( l_43 [393] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2213]    = ( l_43 [394] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2214]    = ( l_43 [395] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2215]    = ( l_43 [396] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2216]    = ( l_43 [397] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2217]    = ( l_43 [398] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[2218]    = ( l_43 [391] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2219]    = ( l_43 [392] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2220]    = ( l_43 [393] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2221]    = ( l_43 [394] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2222]    = ( l_43 [395] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2223]    = ( l_43 [396] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2224]    = ( l_43 [397] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2225]    = ( l_43 [398] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[2226]    = ( l_43 [391] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2227]    = ( l_43 [392] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2228]    = ( l_43 [393] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2229]    = ( l_43 [394] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2230]    = ( l_43 [395] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2231]    = ( l_43 [396] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2232]    = ( l_43 [397] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2233]    = ( l_43 [398] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[2234]    = ( l_43 [391] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2235]    = ( l_43 [392] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2236]    = ( l_43 [393] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2237]    = ( l_43 [394] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2238]    = ( l_43 [395] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2239]    = ( l_43 [396] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2240]    = ( l_43 [397] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2241]    = ( l_43 [398] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[2242]    = ( l_43 [391] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2243]    = ( l_43 [392] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2244]    = ( l_43 [393] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2245]    = ( l_43 [394] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2246]    = ( l_43 [395] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2247]    = ( l_43 [396] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2248]    = ( l_43 [397] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2249]    = ( l_43 [398] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[2250]    = ( l_43 [391] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2251]    = ( l_43 [392] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2252]    = ( l_43 [393] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2253]    = ( l_43 [394] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2254]    = ( l_43 [395] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2255]    = ( l_43 [396] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2256]    = ( l_43 [397] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2257]    = ( l_43 [398] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[2258]    = ( l_43 [391] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2259]    = ( l_43 [392] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2260]    = ( l_43 [393] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2261]    = ( l_43 [394] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2262]    = ( l_43 [395] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2263]    = ( l_43 [396] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2264]    = ( l_43 [397] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2265]    = ( l_43 [398] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[2266]    = ( l_43 [391] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2267]    = ( l_43 [392] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2268]    = ( l_43 [393] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2269]    = ( l_43 [394] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2270]    = ( l_43 [395] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2271]    = ( l_43 [396] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2272]    = ( l_43 [397] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2273]    = ( l_43 [398] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[2274]    = ( l_43 [391] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2275]    = ( l_43 [392] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2276]    = ( l_43 [393] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2277]    = ( l_43 [394] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2278]    = ( l_43 [395] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2279]    = ( l_43 [396] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2280]    = ( l_43 [397] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2281]    = ( l_43 [398] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[2282]    = ( l_43 [391] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2283]    = ( l_43 [392] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2284]    = ( l_43 [393] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2285]    = ( l_43 [394] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2286]    = ( l_43 [395] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2287]    = ( l_43 [396] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2288]    = ( l_43 [397] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2289]    = ( l_43 [398] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[2290]    = ( l_43 [391] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2291]    = ( l_43 [392] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2292]    = ( l_43 [393] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2293]    = ( l_43 [394] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2294]    = ( l_43 [395] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2295]    = ( l_43 [396] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2296]    = ( l_43 [397] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2297]    = ( l_43 [398] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[2298]    = ( l_43 [391] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2299]    = ( l_43 [392] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2300]    = ( l_43 [393] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2301]    = ( l_43 [394] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2302]    = ( l_43 [395] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2303]    = ( l_43 [396] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2304]    = ( l_43 [397] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2305]    = ( l_43 [398] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[2306]    = ( l_43 [391] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2307]    = ( l_43 [392] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2308]    = ( l_43 [393] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2309]    = ( l_43 [394] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2310]    = ( l_43 [395] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2311]    = ( l_43 [396] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2312]    = ( l_43 [397] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2313]    = ( l_43 [398] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[2314]    = ( l_43 [391] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2315]    = ( l_43 [392] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2316]    = ( l_43 [393] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2317]    = ( l_43 [394] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2318]    = ( l_43 [395] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2319]    = ( l_43 [396] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2320]    = ( l_43 [397] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2321]    = ( l_43 [398] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[2322]    = ( l_43 [391] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2323]    = ( l_43 [392] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2324]    = ( l_43 [393] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2325]    = ( l_43 [394] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2326]    = ( l_43 [395] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2327]    = ( l_43 [396] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2328]    = ( l_43 [397] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2329]    = ( l_43 [398] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[2330]    = ( l_43 [391] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2331]    = ( l_43 [392] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2332]    = ( l_43 [393] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2333]    = ( l_43 [394] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2334]    = ( l_43 [395] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2335]    = ( l_43 [396] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2336]    = ( l_43 [397] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2337]    = ( l_43 [398] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[2338]    = ( l_43 [391] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2339]    = ( l_43 [392] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2340]    = ( l_43 [393] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2341]    = ( l_43 [394] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2342]    = ( l_43 [395] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2343]    = ( l_43 [396] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2344]    = ( l_43 [397] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2345]    = ( l_43 [398] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[2346]    = ( l_43 [391] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2347]    = ( l_43 [392] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2348]    = ( l_43 [393] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2349]    = ( l_43 [394] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2350]    = ( l_43 [395] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2351]    = ( l_43 [396] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2352]    = ( l_43 [397] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2353]    = ( l_43 [398] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[2354]    = ( l_43 [391] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2355]    = ( l_43 [392] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2356]    = ( l_43 [393] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2357]    = ( l_43 [394] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2358]    = ( l_43 [395] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2359]    = ( l_43 [396] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2360]    = ( l_43 [397] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2361]    = ( l_43 [398] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[2362]    = ( l_43 [391] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2363]    = ( l_43 [392] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2364]    = ( l_43 [393] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2365]    = ( l_43 [394] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2366]    = ( l_43 [395] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2367]    = ( l_43 [396] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2368]    = ( l_43 [397] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2369]    = ( l_43 [398] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[2370]    = ( l_43 [391] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2371]    = ( l_43 [392] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2372]    = ( l_43 [393] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2373]    = ( l_43 [394] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2374]    = ( l_43 [395] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2375]    = ( l_43 [396] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2376]    = ( l_43 [397] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2377]    = ( l_43 [398] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[2378]    = ( l_43 [391] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2379]    = ( l_43 [392] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2380]    = ( l_43 [393] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2381]    = ( l_43 [394] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2382]    = ( l_43 [395] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2383]    = ( l_43 [396] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2384]    = ( l_43 [397] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2385]    = ( l_43 [398] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[2386]    = ( l_43 [391] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2387]    = ( l_43 [392] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2388]    = ( l_43 [393] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2389]    = ( l_43 [394] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2390]    = ( l_43 [395] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2391]    = ( l_43 [396] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2392]    = ( l_43 [397] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2393]    = ( l_43 [398] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[2394]    = ( l_43 [391] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2395]    = ( l_43 [392] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2396]    = ( l_43 [393] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2397]    = ( l_43 [394] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2398]    = ( l_43 [395] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2399]    = ( l_43 [396] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2400]    = ( l_43 [397] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2401]    = ( l_43 [398] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[2402]    = ( l_43 [391] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2403]    = ( l_43 [392] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2404]    = ( l_43 [393] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2405]    = ( l_43 [394] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2406]    = ( l_43 [395] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2407]    = ( l_43 [396] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2408]    = ( l_43 [397] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2409]    = ( l_43 [398] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[2410]    = ( l_43 [391] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2411]    = ( l_43 [392] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2412]    = ( l_43 [393] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2413]    = ( l_43 [394] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2414]    = ( l_43 [395] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2415]    = ( l_43 [396] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2416]    = ( l_43 [397] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2417]    = ( l_43 [398] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[2418]    = ( l_43 [391] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2419]    = ( l_43 [392] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2420]    = ( l_43 [393] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2421]    = ( l_43 [394] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2422]    = ( l_43 [395] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2423]    = ( l_43 [396] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2424]    = ( l_43 [397] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2425]    = ( l_43 [398] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[2426]    = ( l_43 [391] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2427]    = ( l_43 [392] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2428]    = ( l_43 [393] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2429]    = ( l_43 [394] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2430]    = ( l_43 [395] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2431]    = ( l_43 [396] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2432]    = ( l_43 [397] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2433]    = ( l_43 [398] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[2434]    = ( l_43 [391] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2435]    = ( l_43 [392] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2436]    = ( l_43 [393] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2437]    = ( l_43 [394] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2438]    = ( l_43 [395] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2439]    = ( l_43 [396] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2440]    = ( l_43 [397] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2441]    = ( l_43 [398] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[2442]    = ( l_43 [391] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2443]    = ( l_43 [392] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2444]    = ( l_43 [393] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2445]    = ( l_43 [394] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2446]    = ( l_43 [395] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2447]    = ( l_43 [396] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2448]    = ( l_43 [397] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2449]    = ( l_43 [398] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[2450]    = ( l_43 [391] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2451]    = ( l_43 [392] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2452]    = ( l_43 [393] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2453]    = ( l_43 [394] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2454]    = ( l_43 [395] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2455]    = ( l_43 [396] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2456]    = ( l_43 [397] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2457]    = ( l_43 [398] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[2458]    = ( l_43 [391] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2459]    = ( l_43 [392] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2460]    = ( l_43 [393] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2461]    = ( l_43 [394] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2462]    = ( l_43 [395] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2463]    = ( l_43 [396] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2464]    = ( l_43 [397] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2465]    = ( l_43 [398] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[2466]    = ( l_43 [391] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2467]    = ( l_43 [392] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2468]    = ( l_43 [393] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2469]    = ( l_43 [394] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2470]    = ( l_43 [395] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2471]    = ( l_43 [396] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2472]    = ( l_43 [397] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2473]    = ( l_43 [398] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[2474]    = ( l_43 [391] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2475]    = ( l_43 [392] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2476]    = ( l_43 [393] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2477]    = ( l_43 [394] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2478]    = ( l_43 [395] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2479]    = ( l_43 [396] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2480]    = ( l_43 [397] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2481]    = ( l_43 [398] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[2482]    = ( l_43 [391] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2483]    = ( l_43 [392] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2484]    = ( l_43 [393] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2485]    = ( l_43 [394] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2486]    = ( l_43 [395] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2487]    = ( l_43 [396] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2488]    = ( l_43 [397] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2489]    = ( l_43 [398] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[2490]    = ( l_43 [391] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2491]    = ( l_43 [392] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2492]    = ( l_43 [393] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2493]    = ( l_43 [394] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2494]    = ( l_43 [395] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2495]    = ( l_43 [396] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2496]    = ( l_43 [397] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2497]    = ( l_43 [398] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[2498]    = ( l_43 [391] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2499]    = ( l_43 [392] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2500]    = ( l_43 [393] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2501]    = ( l_43 [394] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2502]    = ( l_43 [395] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2503]    = ( l_43 [396] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2504]    = ( l_43 [397] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2505]    = ( l_43 [398] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[2506]    = ( l_43 [391] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2507]    = ( l_43 [392] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2508]    = ( l_43 [393] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2509]    = ( l_43 [394] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2510]    = ( l_43 [395] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2511]    = ( l_43 [396] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2512]    = ( l_43 [397] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2513]    = ( l_43 [398] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[2514]    = ( l_43 [391] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2515]    = ( l_43 [392] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2516]    = ( l_43 [393] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2517]    = ( l_43 [394] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2518]    = ( l_43 [395] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2519]    = ( l_43 [396] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2520]    = ( l_43 [397] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2521]    = ( l_43 [398] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[2522]    = ( l_43 [391] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2523]    = ( l_43 [392] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2524]    = ( l_43 [393] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2525]    = ( l_43 [394] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2526]    = ( l_43 [395] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2527]    = ( l_43 [396] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2528]    = ( l_43 [397] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2529]    = ( l_43 [398] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[2530]    = ( l_43 [391] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2531]    = ( l_43 [392] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2532]    = ( l_43 [393] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2533]    = ( l_43 [394] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2534]    = ( l_43 [395] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2535]    = ( l_43 [396] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2536]    = ( l_43 [397] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2537]    = ( l_43 [398] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[2538]    = ( l_43 [391] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2539]    = ( l_43 [392] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2540]    = ( l_43 [393] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2541]    = ( l_43 [394] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2542]    = ( l_43 [395] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2543]    = ( l_43 [396] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2544]    = ( l_43 [397] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2545]    = ( l_43 [398] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[2546]    = ( l_43 [391] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2547]    = ( l_43 [392] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2548]    = ( l_43 [393] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2549]    = ( l_43 [394] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2550]    = ( l_43 [395] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2551]    = ( l_43 [396] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2552]    = ( l_43 [397] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2553]    = ( l_43 [398] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[2554]    = ( l_43 [391] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2555]    = ( l_43 [392] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2556]    = ( l_43 [393] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2557]    = ( l_43 [394] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2558]    = ( l_43 [395] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2559]    = ( l_43 [396] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2560]    = ( l_43 [397] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2561]    = ( l_43 [398] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[2562]    = ( l_43 [391] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2563]    = ( l_43 [392] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2564]    = ( l_43 [393] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2565]    = ( l_43 [394] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2566]    = ( l_43 [395] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2567]    = ( l_43 [396] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2568]    = ( l_43 [397] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2569]    = ( l_43 [398] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[2570]    = ( l_43 [391] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2571]    = ( l_43 [392] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2572]    = ( l_43 [393] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2573]    = ( l_43 [394] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2574]    = ( l_43 [395] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2575]    = ( l_43 [396] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2576]    = ( l_43 [397] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2577]    = ( l_43 [398] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[2578]    = ( l_43 [391] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2579]    = ( l_43 [392] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2580]    = ( l_43 [393] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2581]    = ( l_43 [394] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2582]    = ( l_43 [395] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2583]    = ( l_43 [396] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2584]    = ( l_43 [397] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2585]    = ( l_43 [398] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[2586]    = ( l_43 [391] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2587]    = ( l_43 [392] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2588]    = ( l_43 [393] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2589]    = ( l_43 [394] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2590]    = ( l_43 [395] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2591]    = ( l_43 [396] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2592]    = ( l_43 [397] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2593]    = ( l_43 [398] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[2594]    = ( l_43 [391] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2595]    = ( l_43 [392] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2596]    = ( l_43 [393] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2597]    = ( l_43 [394] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2598]    = ( l_43 [395] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2599]    = ( l_43 [396] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2600]    = ( l_43 [397] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2601]    = ( l_43 [398] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[2602]    = ( l_43 [391] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2603]    = ( l_43 [392] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2604]    = ( l_43 [393] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2605]    = ( l_43 [394] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2606]    = ( l_43 [395] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2607]    = ( l_43 [396] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2608]    = ( l_43 [397] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2609]    = ( l_43 [398] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[2610]    = ( l_43 [391] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2611]    = ( l_43 [392] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2612]    = ( l_43 [393] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2613]    = ( l_43 [394] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2614]    = ( l_43 [395] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2615]    = ( l_43 [396] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2616]    = ( l_43 [397] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2617]    = ( l_43 [398] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[2618]    = ( l_43 [391] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2619]    = ( l_43 [392] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2620]    = ( l_43 [393] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2621]    = ( l_43 [394] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2622]    = ( l_43 [395] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2623]    = ( l_43 [396] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2624]    = ( l_43 [397] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2625]    = ( l_43 [398] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[2626]    = ( l_43 [391] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2627]    = ( l_43 [392] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2628]    = ( l_43 [393] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2629]    = ( l_43 [394] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2630]    = ( l_43 [395] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2631]    = ( l_43 [396] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2632]    = ( l_43 [397] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2633]    = ( l_43 [398] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[2634]    = ( l_43 [391] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2635]    = ( l_43 [392] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2636]    = ( l_43 [393] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2637]    = ( l_43 [394] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2638]    = ( l_43 [395] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2639]    = ( l_43 [396] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2640]    = ( l_43 [397] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2641]    = ( l_43 [398] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[2642]    = ( l_43 [391] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2643]    = ( l_43 [392] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2644]    = ( l_43 [393] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2645]    = ( l_43 [394] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2646]    = ( l_43 [395] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2647]    = ( l_43 [396] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2648]    = ( l_43 [397] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2649]    = ( l_43 [398] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[2650]    = ( l_43 [391] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2651]    = ( l_43 [392] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2652]    = ( l_43 [393] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2653]    = ( l_43 [394] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2654]    = ( l_43 [395] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2655]    = ( l_43 [396] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2656]    = ( l_43 [397] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2657]    = ( l_43 [398] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[2658]    = ( l_43 [391] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2659]    = ( l_43 [392] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2660]    = ( l_43 [393] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2661]    = ( l_43 [394] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2662]    = ( l_43 [395] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2663]    = ( l_43 [396] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2664]    = ( l_43 [397] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2665]    = ( l_43 [398] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[2666]    = ( l_43 [391] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2667]    = ( l_43 [392] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2668]    = ( l_43 [393] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2669]    = ( l_43 [394] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2670]    = ( l_43 [395] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2671]    = ( l_43 [396] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2672]    = ( l_43 [397] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2673]    = ( l_43 [398] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[2674]    = ( l_43 [391] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2675]    = ( l_43 [392] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2676]    = ( l_43 [393] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2677]    = ( l_43 [394] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2678]    = ( l_43 [395] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2679]    = ( l_43 [396] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2680]    = ( l_43 [397] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2681]    = ( l_43 [398] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[2682]    = ( l_43 [391] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2683]    = ( l_43 [392] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2684]    = ( l_43 [393] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2685]    = ( l_43 [394] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2686]    = ( l_43 [395] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2687]    = ( l_43 [396] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2688]    = ( l_43 [397] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2689]    = ( l_43 [398] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[2690]    = ( l_43 [391] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2691]    = ( l_43 [392] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2692]    = ( l_43 [393] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2693]    = ( l_43 [394] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2694]    = ( l_43 [395] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2695]    = ( l_43 [396] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2696]    = ( l_43 [397] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2697]    = ( l_43 [398] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[2698]    = ( l_43 [391] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2699]    = ( l_43 [392] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2700]    = ( l_43 [393] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2701]    = ( l_43 [394] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2702]    = ( l_43 [395] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2703]    = ( l_43 [396] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2704]    = ( l_43 [397] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2705]    = ( l_43 [398] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[2706]    = ( l_43 [391] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2707]    = ( l_43 [392] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2708]    = ( l_43 [393] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2709]    = ( l_43 [394] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2710]    = ( l_43 [395] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2711]    = ( l_43 [396] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2712]    = ( l_43 [397] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2713]    = ( l_43 [398] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[2714]    = ( l_43 [391] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2715]    = ( l_43 [392] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2716]    = ( l_43 [393] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2717]    = ( l_43 [394] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2718]    = ( l_43 [395] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2719]    = ( l_43 [396] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2720]    = ( l_43 [397] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2721]    = ( l_43 [398] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[2722]    = ( l_43 [391] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2723]    = ( l_43 [392] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2724]    = ( l_43 [393] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2725]    = ( l_43 [394] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2726]    = ( l_43 [395] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2727]    = ( l_43 [396] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2728]    = ( l_43 [397] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2729]    = ( l_43 [398] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[2730]    = ( l_43 [391] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2731]    = ( l_43 [392] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2732]    = ( l_43 [393] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2733]    = ( l_43 [394] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2734]    = ( l_43 [395] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2735]    = ( l_43 [396] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2736]    = ( l_43 [397] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2737]    = ( l_43 [398] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[2738]    = ( l_43 [391] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2739]    = ( l_43 [392] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2740]    = ( l_43 [393] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2741]    = ( l_43 [394] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2742]    = ( l_43 [395] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2743]    = ( l_43 [396] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2744]    = ( l_43 [397] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2745]    = ( l_43 [398] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[2746]    = ( l_43 [391] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2747]    = ( l_43 [392] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2748]    = ( l_43 [393] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2749]    = ( l_43 [394] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2750]    = ( l_43 [395] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2751]    = ( l_43 [396] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2752]    = ( l_43 [397] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2753]    = ( l_43 [398] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[2754]    = ( l_43 [391] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2755]    = ( l_43 [392] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2756]    = ( l_43 [393] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2757]    = ( l_43 [394] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2758]    = ( l_43 [395] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2759]    = ( l_43 [396] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2760]    = ( l_43 [397] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2761]    = ( l_43 [398] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[2762]    = ( l_43 [391] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2763]    = ( l_43 [392] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2764]    = ( l_43 [393] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2765]    = ( l_43 [394] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2766]    = ( l_43 [395] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2767]    = ( l_43 [396] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2768]    = ( l_43 [397] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2769]    = ( l_43 [398] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[2770]    = ( l_43 [391] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2771]    = ( l_43 [392] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2772]    = ( l_43 [393] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2773]    = ( l_43 [394] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2774]    = ( l_43 [395] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2775]    = ( l_43 [396] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2776]    = ( l_43 [397] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2777]    = ( l_43 [398] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[2778]    = ( l_43 [391] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2779]    = ( l_43 [392] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2780]    = ( l_43 [393] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2781]    = ( l_43 [394] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2782]    = ( l_43 [395] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2783]    = ( l_43 [396] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2784]    = ( l_43 [397] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2785]    = ( l_43 [398] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[2786]    = ( l_43 [391] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2787]    = ( l_43 [392] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2788]    = ( l_43 [393] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2789]    = ( l_43 [394] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2790]    = ( l_43 [395] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2791]    = ( l_43 [396] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2792]    = ( l_43 [397] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2793]    = ( l_43 [398] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[2794]    = ( l_43 [391] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2795]    = ( l_43 [392] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2796]    = ( l_43 [393] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2797]    = ( l_43 [394] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2798]    = ( l_43 [395] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2799]    = ( l_43 [396] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2800]    = ( l_43 [397] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2801]    = ( l_43 [398] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[2802]    = ( l_43 [391] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2803]    = ( l_43 [392] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2804]    = ( l_43 [393] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2805]    = ( l_43 [394] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2806]    = ( l_43 [395] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2807]    = ( l_43 [396] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2808]    = ( l_43 [397] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2809]    = ( l_43 [398] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[2810]    = ( l_43 [391] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2811]    = ( l_43 [392] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2812]    = ( l_43 [393] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2813]    = ( l_43 [394] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2814]    = ( l_43 [395] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2815]    = ( l_43 [396] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2816]    = ( l_43 [397] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2817]    = ( l_43 [398] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[2818]    = ( l_43 [391] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2819]    = ( l_43 [392] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2820]    = ( l_43 [393] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2821]    = ( l_43 [394] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2822]    = ( l_43 [395] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2823]    = ( l_43 [396] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2824]    = ( l_43 [397] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2825]    = ( l_43 [398] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[2826]    = ( l_43 [391] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2827]    = ( l_43 [392] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2828]    = ( l_43 [393] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2829]    = ( l_43 [394] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2830]    = ( l_43 [395] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2831]    = ( l_43 [396] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2832]    = ( l_43 [397] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2833]    = ( l_43 [398] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[2834]    = ( l_43 [391] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2835]    = ( l_43 [392] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2836]    = ( l_43 [393] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2837]    = ( l_43 [394] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2838]    = ( l_43 [395] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2839]    = ( l_43 [396] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2840]    = ( l_43 [397] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2841]    = ( l_43 [398] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[2842]    = ( l_43 [391] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2843]    = ( l_43 [392] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2844]    = ( l_43 [393] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2845]    = ( l_43 [394] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2846]    = ( l_43 [395] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2847]    = ( l_43 [396] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2848]    = ( l_43 [397] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2849]    = ( l_43 [398] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[2850]    = ( l_43 [391] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2851]    = ( l_43 [392] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2852]    = ( l_43 [393] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2853]    = ( l_43 [394] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2854]    = ( l_43 [395] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2855]    = ( l_43 [396] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2856]    = ( l_43 [397] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2857]    = ( l_43 [398] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[2858]    = ( l_43 [391] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2859]    = ( l_43 [392] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2860]    = ( l_43 [393] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2861]    = ( l_43 [394] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2862]    = ( l_43 [395] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2863]    = ( l_43 [396] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2864]    = ( l_43 [397] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2865]    = ( l_43 [398] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[2866]    = ( l_43 [391] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2867]    = ( l_43 [392] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2868]    = ( l_43 [393] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2869]    = ( l_43 [394] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2870]    = ( l_43 [395] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2871]    = ( l_43 [396] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2872]    = ( l_43 [397] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2873]    = ( l_43 [398] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[2874]    = ( l_43 [391] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2875]    = ( l_43 [392] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2876]    = ( l_43 [393] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2877]    = ( l_43 [394] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2878]    = ( l_43 [395] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2879]    = ( l_43 [396] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2880]    = ( l_43 [397] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2881]    = ( l_43 [398] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[2882]    = ( l_43 [391] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2883]    = ( l_43 [392] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2884]    = ( l_43 [393] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2885]    = ( l_43 [394] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2886]    = ( l_43 [395] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2887]    = ( l_43 [396] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2888]    = ( l_43 [397] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2889]    = ( l_43 [398] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[2890]    = ( l_43 [391] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2891]    = ( l_43 [392] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2892]    = ( l_43 [393] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2893]    = ( l_43 [394] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2894]    = ( l_43 [395] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2895]    = ( l_43 [396] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2896]    = ( l_43 [397] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2897]    = ( l_43 [398] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[2898]    = ( l_43 [391] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2899]    = ( l_43 [392] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2900]    = ( l_43 [393] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2901]    = ( l_43 [394] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2902]    = ( l_43 [395] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2903]    = ( l_43 [396] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2904]    = ( l_43 [397] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2905]    = ( l_43 [398] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[2906]    = ( l_43 [391] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2907]    = ( l_43 [392] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2908]    = ( l_43 [393] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2909]    = ( l_43 [394] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2910]    = ( l_43 [395] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2911]    = ( l_43 [396] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2912]    = ( l_43 [397] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2913]    = ( l_43 [398] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[2914]    = ( l_43 [391] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2915]    = ( l_43 [392] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2916]    = ( l_43 [393] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2917]    = ( l_43 [394] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2918]    = ( l_43 [395] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2919]    = ( l_43 [396] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2920]    = ( l_43 [397] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2921]    = ( l_43 [398] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[2922]    = ( l_43 [391] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2923]    = ( l_43 [392] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2924]    = ( l_43 [393] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2925]    = ( l_43 [394] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2926]    = ( l_43 [395] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2927]    = ( l_43 [396] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2928]    = ( l_43 [397] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2929]    = ( l_43 [398] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[2930]    = ( l_43 [391] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2931]    = ( l_43 [392] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2932]    = ( l_43 [393] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2933]    = ( l_43 [394] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2934]    = ( l_43 [395] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2935]    = ( l_43 [396] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2936]    = ( l_43 [397] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2937]    = ( l_43 [398] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[2938]    = ( l_43 [391] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2939]    = ( l_43 [392] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2940]    = ( l_43 [393] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2941]    = ( l_43 [394] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2942]    = ( l_43 [395] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2943]    = ( l_43 [396] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2944]    = ( l_43 [397] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2945]    = ( l_43 [398] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[2946]    = ( l_43 [391] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2947]    = ( l_43 [392] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2948]    = ( l_43 [393] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2949]    = ( l_43 [394] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2950]    = ( l_43 [395] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2951]    = ( l_43 [396] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2952]    = ( l_43 [397] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2953]    = ( l_43 [398] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[2954]    = ( l_43 [391] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2955]    = ( l_43 [392] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2956]    = ( l_43 [393] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2957]    = ( l_43 [394] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2958]    = ( l_43 [395] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2959]    = ( l_43 [396] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2960]    = ( l_43 [397] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2961]    = ( l_43 [398] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[2962]    = ( l_43 [391] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2963]    = ( l_43 [392] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2964]    = ( l_43 [393] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2965]    = ( l_43 [394] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2966]    = ( l_43 [395] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2967]    = ( l_43 [396] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2968]    = ( l_43 [397] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2969]    = ( l_43 [398] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[2970]    = ( l_43 [391] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2971]    = ( l_43 [392] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2972]    = ( l_43 [393] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2973]    = ( l_43 [394] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2974]    = ( l_43 [395] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2975]    = ( l_43 [396] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2976]    = ( l_43 [397] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2977]    = ( l_43 [398] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[2978]    = ( l_43 [391] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2979]    = ( l_43 [392] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2980]    = ( l_43 [393] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2981]    = ( l_43 [394] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2982]    = ( l_43 [395] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2983]    = ( l_43 [396] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2984]    = ( l_43 [397] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2985]    = ( l_43 [398] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[2986]    = ( l_43 [391] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2987]    = ( l_43 [392] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2988]    = ( l_43 [393] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2989]    = ( l_43 [394] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2990]    = ( l_43 [395] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2991]    = ( l_43 [396] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2992]    = ( l_43 [397] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2993]    = ( l_43 [398] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[2994]    = ( l_43 [391] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[2995]    = ( l_43 [392] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[2996]    = ( l_43 [393] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[2997]    = ( l_43 [394] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[2998]    = ( l_43 [395] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[2999]    = ( l_43 [396] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[3000]    = ( l_43 [397] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[3001]    = ( l_43 [398] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[3002]    = ( l_43 [391] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3003]    = ( l_43 [392] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3004]    = ( l_43 [393] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3005]    = ( l_43 [394] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3006]    = ( l_43 [395] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3007]    = ( l_43 [396] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3008]    = ( l_43 [397] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3009]    = ( l_43 [398] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[3010]    = ( l_43 [391] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3011]    = ( l_43 [392] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3012]    = ( l_43 [393] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3013]    = ( l_43 [394] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3014]    = ( l_43 [395] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3015]    = ( l_43 [396] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3016]    = ( l_43 [397] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3017]    = ( l_43 [398] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[3018]    = ( l_43 [391] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3019]    = ( l_43 [392] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3020]    = ( l_43 [393] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3021]    = ( l_43 [394] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3022]    = ( l_43 [395] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3023]    = ( l_43 [396] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3024]    = ( l_43 [397] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3025]    = ( l_43 [398] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[3026]    = ( l_43 [391] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3027]    = ( l_43 [392] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3028]    = ( l_43 [393] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3029]    = ( l_43 [394] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3030]    = ( l_43 [395] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3031]    = ( l_43 [396] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3032]    = ( l_43 [397] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3033]    = ( l_43 [398] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[3034]    = ( l_43 [391] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3035]    = ( l_43 [392] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3036]    = ( l_43 [393] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3037]    = ( l_43 [394] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3038]    = ( l_43 [395] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3039]    = ( l_43 [396] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3040]    = ( l_43 [397] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3041]    = ( l_43 [398] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[3042]    = ( l_43 [391] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3043]    = ( l_43 [392] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3044]    = ( l_43 [393] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3045]    = ( l_43 [394] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3046]    = ( l_43 [395] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3047]    = ( l_43 [396] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3048]    = ( l_43 [397] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3049]    = ( l_43 [398] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[3050]    = ( l_43 [391] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3051]    = ( l_43 [392] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3052]    = ( l_43 [393] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3053]    = ( l_43 [394] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3054]    = ( l_43 [395] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3055]    = ( l_43 [396] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3056]    = ( l_43 [397] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3057]    = ( l_43 [398] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[3058]    = ( l_43 [391] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3059]    = ( l_43 [392] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3060]    = ( l_43 [393] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3061]    = ( l_43 [394] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3062]    = ( l_43 [395] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3063]    = ( l_43 [396] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3064]    = ( l_43 [397] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3065]    = ( l_43 [398] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[3066]    = ( l_43 [391] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3067]    = ( l_43 [392] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3068]    = ( l_43 [393] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3069]    = ( l_43 [394] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3070]    = ( l_43 [395] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3071]    = ( l_43 [396] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3072]    = ( l_43 [397] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3073]    = ( l_43 [398] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[3074]    = ( l_43 [391] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3075]    = ( l_43 [392] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3076]    = ( l_43 [393] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3077]    = ( l_43 [394] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3078]    = ( l_43 [395] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3079]    = ( l_43 [396] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3080]    = ( l_43 [397] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3081]    = ( l_43 [398] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[3082]    = ( l_43 [391] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3083]    = ( l_43 [392] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3084]    = ( l_43 [393] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3085]    = ( l_43 [394] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3086]    = ( l_43 [395] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3087]    = ( l_43 [396] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3088]    = ( l_43 [397] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3089]    = ( l_43 [398] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[3090]    = ( l_43 [391] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3091]    = ( l_43 [392] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3092]    = ( l_43 [393] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3093]    = ( l_43 [394] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3094]    = ( l_43 [395] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3095]    = ( l_43 [396] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3096]    = ( l_43 [397] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3097]    = ( l_43 [398] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[3098]    = ( l_43 [391] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3099]    = ( l_43 [392] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3100]    = ( l_43 [393] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3101]    = ( l_43 [394] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3102]    = ( l_43 [395] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3103]    = ( l_43 [396] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3104]    = ( l_43 [397] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3105]    = ( l_43 [398] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[3106]    = ( l_43 [391] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3107]    = ( l_43 [392] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3108]    = ( l_43 [393] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3109]    = ( l_43 [394] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3110]    = ( l_43 [395] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3111]    = ( l_43 [396] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3112]    = ( l_43 [397] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3113]    = ( l_43 [398] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[3114]    = ( l_43 [391] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3115]    = ( l_43 [392] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3116]    = ( l_43 [393] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3117]    = ( l_43 [394] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3118]    = ( l_43 [395] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3119]    = ( l_43 [396] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3120]    = ( l_43 [397] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3121]    = ( l_43 [398] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[3122]    = ( l_43 [391] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3123]    = ( l_43 [392] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3124]    = ( l_43 [393] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3125]    = ( l_43 [394] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3126]    = ( l_43 [395] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3127]    = ( l_43 [396] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3128]    = ( l_43 [397] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3129]    = ( l_43 [398] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[3130]    = ( l_43 [391] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3131]    = ( l_43 [392] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3132]    = ( l_43 [393] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3133]    = ( l_43 [394] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3134]    = ( l_43 [395] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3135]    = ( l_43 [396] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3136]    = ( l_43 [397] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3137]    = ( l_43 [398] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[3138]    = ( l_43 [391] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3139]    = ( l_43 [392] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3140]    = ( l_43 [393] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3141]    = ( l_43 [394] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3142]    = ( l_43 [395] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3143]    = ( l_43 [396] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3144]    = ( l_43 [397] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3145]    = ( l_43 [398] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[3146]    = ( l_43 [391] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3147]    = ( l_43 [392] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3148]    = ( l_43 [393] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3149]    = ( l_43 [394] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3150]    = ( l_43 [395] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3151]    = ( l_43 [396] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3152]    = ( l_43 [397] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3153]    = ( l_43 [398] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[3154]    = ( l_43 [391] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3155]    = ( l_43 [392] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3156]    = ( l_43 [393] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3157]    = ( l_43 [394] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3158]    = ( l_43 [395] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3159]    = ( l_43 [396] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3160]    = ( l_43 [397] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3161]    = ( l_43 [398] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[3162]    = ( l_43 [391] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3163]    = ( l_43 [392] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3164]    = ( l_43 [393] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3165]    = ( l_43 [394] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3166]    = ( l_43 [395] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3167]    = ( l_43 [396] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3168]    = ( l_43 [397] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3169]    = ( l_43 [398] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[3170]    = ( l_43 [391] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3171]    = ( l_43 [392] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3172]    = ( l_43 [393] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3173]    = ( l_43 [394] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3174]    = ( l_43 [395] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3175]    = ( l_43 [396] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3176]    = ( l_43 [397] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3177]    = ( l_43 [398] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[3178]    = ( l_43 [391] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3179]    = ( l_43 [392] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3180]    = ( l_43 [393] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3181]    = ( l_43 [394] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3182]    = ( l_43 [395] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3183]    = ( l_43 [396] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3184]    = ( l_43 [397] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3185]    = ( l_43 [398] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[3186]    = ( l_43 [391] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3187]    = ( l_43 [392] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3188]    = ( l_43 [393] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3189]    = ( l_43 [394] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3190]    = ( l_43 [395] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3191]    = ( l_43 [396] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3192]    = ( l_43 [397] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3193]    = ( l_43 [398] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[3194]    = ( l_43 [391] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3195]    = ( l_43 [392] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3196]    = ( l_43 [393] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3197]    = ( l_43 [394] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3198]    = ( l_43 [395] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3199]    = ( l_43 [396] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3200]    = ( l_43 [397] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3201]    = ( l_43 [398] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[3202]    = ( l_43 [391] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3203]    = ( l_43 [392] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3204]    = ( l_43 [393] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3205]    = ( l_43 [394] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3206]    = ( l_43 [395] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3207]    = ( l_43 [396] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3208]    = ( l_43 [397] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3209]    = ( l_43 [398] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[3210]    = ( l_43 [391] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3211]    = ( l_43 [392] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3212]    = ( l_43 [393] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3213]    = ( l_43 [394] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3214]    = ( l_43 [395] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3215]    = ( l_43 [396] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3216]    = ( l_43 [397] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3217]    = ( l_43 [398] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[3218]    = ( l_43 [391] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3219]    = ( l_43 [392] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3220]    = ( l_43 [393] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3221]    = ( l_43 [394] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3222]    = ( l_43 [395] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3223]    = ( l_43 [396] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3224]    = ( l_43 [397] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3225]    = ( l_43 [398] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[3226]    = ( l_43 [391] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3227]    = ( l_43 [392] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3228]    = ( l_43 [393] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3229]    = ( l_43 [394] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3230]    = ( l_43 [395] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3231]    = ( l_43 [396] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3232]    = ( l_43 [397] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3233]    = ( l_43 [398] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[3234]    = ( l_43 [391] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3235]    = ( l_43 [392] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3236]    = ( l_43 [393] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3237]    = ( l_43 [394] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3238]    = ( l_43 [395] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3239]    = ( l_43 [396] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3240]    = ( l_43 [397] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3241]    = ( l_43 [398] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[3242]    = ( l_43 [391] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3243]    = ( l_43 [392] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3244]    = ( l_43 [393] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3245]    = ( l_43 [394] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3246]    = ( l_43 [395] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3247]    = ( l_43 [396] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3248]    = ( l_43 [397] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3249]    = ( l_43 [398] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[3250]    = ( l_43 [391] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3251]    = ( l_43 [392] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3252]    = ( l_43 [393] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3253]    = ( l_43 [394] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3254]    = ( l_43 [395] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3255]    = ( l_43 [396] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3256]    = ( l_43 [397] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3257]    = ( l_43 [398] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[3258]    = ( l_43 [391] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3259]    = ( l_43 [392] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3260]    = ( l_43 [393] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3261]    = ( l_43 [394] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3262]    = ( l_43 [395] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3263]    = ( l_43 [396] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3264]    = ( l_43 [397] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3265]    = ( l_43 [398] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[3266]    = ( l_43 [391] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3267]    = ( l_43 [392] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3268]    = ( l_43 [393] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3269]    = ( l_43 [394] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3270]    = ( l_43 [395] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3271]    = ( l_43 [396] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3272]    = ( l_43 [397] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3273]    = ( l_43 [398] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[3274]    = ( l_43 [391] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3275]    = ( l_43 [392] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3276]    = ( l_43 [393] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3277]    = ( l_43 [394] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3278]    = ( l_43 [395] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3279]    = ( l_43 [396] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3280]    = ( l_43 [397] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3281]    = ( l_43 [398] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[3282]    = ( l_43 [391] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3283]    = ( l_43 [392] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3284]    = ( l_43 [393] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3285]    = ( l_43 [394] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3286]    = ( l_43 [395] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3287]    = ( l_43 [396] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3288]    = ( l_43 [397] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3289]    = ( l_43 [398] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[3290]    = ( l_43 [391] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3291]    = ( l_43 [392] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3292]    = ( l_43 [393] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3293]    = ( l_43 [394] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3294]    = ( l_43 [395] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3295]    = ( l_43 [396] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3296]    = ( l_43 [397] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3297]    = ( l_43 [398] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[3298]    = ( l_43 [391] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3299]    = ( l_43 [392] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3300]    = ( l_43 [393] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3301]    = ( l_43 [394] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3302]    = ( l_43 [395] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3303]    = ( l_43 [396] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3304]    = ( l_43 [397] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3305]    = ( l_43 [398] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[3306]    = ( l_43 [391] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3307]    = ( l_43 [392] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3308]    = ( l_43 [393] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3309]    = ( l_43 [394] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3310]    = ( l_43 [395] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3311]    = ( l_43 [396] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3312]    = ( l_43 [397] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3313]    = ( l_43 [398] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[3314]    = ( l_43 [391] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3315]    = ( l_43 [392] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3316]    = ( l_43 [393] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3317]    = ( l_43 [394] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3318]    = ( l_43 [395] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3319]    = ( l_43 [396] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3320]    = ( l_43 [397] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3321]    = ( l_43 [398] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[3322]    = ( l_43 [391] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3323]    = ( l_43 [392] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3324]    = ( l_43 [393] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3325]    = ( l_43 [394] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3326]    = ( l_43 [395] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3327]    = ( l_43 [396] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3328]    = ( l_43 [397] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3329]    = ( l_43 [398] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[3330]    = ( l_43 [391] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3331]    = ( l_43 [392] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3332]    = ( l_43 [393] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3333]    = ( l_43 [394] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3334]    = ( l_43 [395] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3335]    = ( l_43 [396] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3336]    = ( l_43 [397] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3337]    = ( l_43 [398] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[3338]    = ( l_43 [391] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3339]    = ( l_43 [392] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3340]    = ( l_43 [393] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3341]    = ( l_43 [394] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3342]    = ( l_43 [395] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3343]    = ( l_43 [396] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3344]    = ( l_43 [397] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3345]    = ( l_43 [398] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[3346]    = ( l_43 [391] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3347]    = ( l_43 [392] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3348]    = ( l_43 [393] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3349]    = ( l_43 [394] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3350]    = ( l_43 [395] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3351]    = ( l_43 [396] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3352]    = ( l_43 [397] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3353]    = ( l_43 [398] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[3354]    = ( l_43 [391] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3355]    = ( l_43 [392] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3356]    = ( l_43 [393] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3357]    = ( l_43 [394] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3358]    = ( l_43 [395] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3359]    = ( l_43 [396] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3360]    = ( l_43 [397] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3361]    = ( l_43 [398] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[3362]    = ( l_43 [391] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3363]    = ( l_43 [392] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3364]    = ( l_43 [393] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3365]    = ( l_43 [394] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3366]    = ( l_43 [395] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3367]    = ( l_43 [396] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3368]    = ( l_43 [397] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3369]    = ( l_43 [398] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[3370]    = ( l_43 [391] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3371]    = ( l_43 [392] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3372]    = ( l_43 [393] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3373]    = ( l_43 [394] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3374]    = ( l_43 [395] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3375]    = ( l_43 [396] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3376]    = ( l_43 [397] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3377]    = ( l_43 [398] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[3378]    = ( l_43 [391] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3379]    = ( l_43 [392] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3380]    = ( l_43 [393] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3381]    = ( l_43 [394] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3382]    = ( l_43 [395] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3383]    = ( l_43 [396] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3384]    = ( l_43 [397] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3385]    = ( l_43 [398] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[3386]    = ( l_43 [391] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3387]    = ( l_43 [392] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3388]    = ( l_43 [393] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3389]    = ( l_43 [394] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3390]    = ( l_43 [395] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3391]    = ( l_43 [396] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3392]    = ( l_43 [397] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3393]    = ( l_43 [398] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[3394]    = ( l_43 [391] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3395]    = ( l_43 [392] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3396]    = ( l_43 [393] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3397]    = ( l_43 [394] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3398]    = ( l_43 [395] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3399]    = ( l_43 [396] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3400]    = ( l_43 [397] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3401]    = ( l_43 [398] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[3402]    = ( l_43 [391] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3403]    = ( l_43 [392] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3404]    = ( l_43 [393] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3405]    = ( l_43 [394] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3406]    = ( l_43 [395] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3407]    = ( l_43 [396] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3408]    = ( l_43 [397] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3409]    = ( l_43 [398] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[3410]    = ( l_43 [391] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3411]    = ( l_43 [392] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3412]    = ( l_43 [393] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3413]    = ( l_43 [394] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3414]    = ( l_43 [395] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3415]    = ( l_43 [396] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3416]    = ( l_43 [397] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3417]    = ( l_43 [398] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[3418]    = ( l_43 [391] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3419]    = ( l_43 [392] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3420]    = ( l_43 [393] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3421]    = ( l_43 [394] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3422]    = ( l_43 [395] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3423]    = ( l_43 [396] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3424]    = ( l_43 [397] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3425]    = ( l_43 [398] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[3426]    = ( l_43 [391] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3427]    = ( l_43 [392] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3428]    = ( l_43 [393] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3429]    = ( l_43 [394] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3430]    = ( l_43 [395] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3431]    = ( l_43 [396] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3432]    = ( l_43 [397] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3433]    = ( l_43 [398] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[3434]    = ( l_43 [391] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3435]    = ( l_43 [392] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3436]    = ( l_43 [393] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3437]    = ( l_43 [394] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3438]    = ( l_43 [395] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3439]    = ( l_43 [396] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3440]    = ( l_43 [397] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3441]    = ( l_43 [398] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[3442]    = ( l_43 [391] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3443]    = ( l_43 [392] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3444]    = ( l_43 [393] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3445]    = ( l_43 [394] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3446]    = ( l_43 [395] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3447]    = ( l_43 [396] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3448]    = ( l_43 [397] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3449]    = ( l_43 [398] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[3450]    = ( l_43 [391] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3451]    = ( l_43 [392] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3452]    = ( l_43 [393] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3453]    = ( l_43 [394] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3454]    = ( l_43 [395] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3455]    = ( l_43 [396] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3456]    = ( l_43 [397] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3457]    = ( l_43 [398] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[3458]    = ( l_43 [391] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3459]    = ( l_43 [392] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3460]    = ( l_43 [393] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3461]    = ( l_43 [394] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3462]    = ( l_43 [395] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3463]    = ( l_43 [396] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3464]    = ( l_43 [397] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3465]    = ( l_43 [398] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[3466]    = ( l_43 [391] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3467]    = ( l_43 [392] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3468]    = ( l_43 [393] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3469]    = ( l_43 [394] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3470]    = ( l_43 [395] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3471]    = ( l_43 [396] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3472]    = ( l_43 [397] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3473]    = ( l_43 [398] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[3474]    = ( l_43 [391] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3475]    = ( l_43 [392] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3476]    = ( l_43 [393] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3477]    = ( l_43 [394] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3478]    = ( l_43 [395] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3479]    = ( l_43 [396] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3480]    = ( l_43 [397] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3481]    = ( l_43 [398] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[3482]    = ( l_43 [391] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3483]    = ( l_43 [392] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3484]    = ( l_43 [393] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3485]    = ( l_43 [394] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3486]    = ( l_43 [395] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3487]    = ( l_43 [396] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3488]    = ( l_43 [397] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3489]    = ( l_43 [398] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[3490]    = ( l_43 [391] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3491]    = ( l_43 [392] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3492]    = ( l_43 [393] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3493]    = ( l_43 [394] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3494]    = ( l_43 [395] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3495]    = ( l_43 [396] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3496]    = ( l_43 [397] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3497]    = ( l_43 [398] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[3498]    = ( l_43 [391] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3499]    = ( l_43 [392] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3500]    = ( l_43 [393] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3501]    = ( l_43 [394] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3502]    = ( l_43 [395] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3503]    = ( l_43 [396] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3504]    = ( l_43 [397] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3505]    = ( l_43 [398] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[3506]    = ( l_43 [391] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3507]    = ( l_43 [392] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3508]    = ( l_43 [393] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3509]    = ( l_43 [394] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3510]    = ( l_43 [395] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3511]    = ( l_43 [396] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3512]    = ( l_43 [397] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3513]    = ( l_43 [398] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[3514]    = ( l_43 [391] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3515]    = ( l_43 [392] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3516]    = ( l_43 [393] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3517]    = ( l_43 [394] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3518]    = ( l_43 [395] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3519]    = ( l_43 [396] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3520]    = ( l_43 [397] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3521]    = ( l_43 [398] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[3522]    = ( l_43 [391] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3523]    = ( l_43 [392] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3524]    = ( l_43 [393] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3525]    = ( l_43 [394] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3526]    = ( l_43 [395] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3527]    = ( l_43 [396] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3528]    = ( l_43 [397] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3529]    = ( l_43 [398] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[3530]    = ( l_43 [391] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3531]    = ( l_43 [392] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3532]    = ( l_43 [393] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3533]    = ( l_43 [394] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3534]    = ( l_43 [395] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3535]    = ( l_43 [396] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3536]    = ( l_43 [397] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3537]    = ( l_43 [398] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[3538]    = ( l_43 [391] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3539]    = ( l_43 [392] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3540]    = ( l_43 [393] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3541]    = ( l_43 [394] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3542]    = ( l_43 [395] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3543]    = ( l_43 [396] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3544]    = ( l_43 [397] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3545]    = ( l_43 [398] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[3546]    = ( l_43 [391] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3547]    = ( l_43 [392] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3548]    = ( l_43 [393] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3549]    = ( l_43 [394] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3550]    = ( l_43 [395] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3551]    = ( l_43 [396] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3552]    = ( l_43 [397] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3553]    = ( l_43 [398] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[3554]    = ( l_43 [391] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3555]    = ( l_43 [392] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3556]    = ( l_43 [393] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3557]    = ( l_43 [394] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3558]    = ( l_43 [395] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3559]    = ( l_43 [396] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3560]    = ( l_43 [397] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3561]    = ( l_43 [398] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[3562]    = ( l_43 [391] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3563]    = ( l_43 [392] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3564]    = ( l_43 [393] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3565]    = ( l_43 [394] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3566]    = ( l_43 [395] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3567]    = ( l_43 [396] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3568]    = ( l_43 [397] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3569]    = ( l_43 [398] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[3570]    = ( l_43 [391] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3571]    = ( l_43 [392] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3572]    = ( l_43 [393] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3573]    = ( l_43 [394] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3574]    = ( l_43 [395] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3575]    = ( l_43 [396] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3576]    = ( l_43 [397] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3577]    = ( l_43 [398] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[3578]    = ( l_43 [391] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3579]    = ( l_43 [392] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3580]    = ( l_43 [393] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3581]    = ( l_43 [394] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3582]    = ( l_43 [395] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3583]    = ( l_43 [396] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3584]    = ( l_43 [397] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3585]    = ( l_43 [398] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[3586]    = ( l_43 [391] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3587]    = ( l_43 [392] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3588]    = ( l_43 [393] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3589]    = ( l_43 [394] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3590]    = ( l_43 [395] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3591]    = ( l_43 [396] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3592]    = ( l_43 [397] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3593]    = ( l_43 [398] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[3594]    = ( l_43 [391] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3595]    = ( l_43 [392] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3596]    = ( l_43 [393] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3597]    = ( l_43 [394] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3598]    = ( l_43 [395] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3599]    = ( l_43 [396] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3600]    = ( l_43 [397] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3601]    = ( l_43 [398] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[3602]    = ( l_43 [391] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3603]    = ( l_43 [392] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3604]    = ( l_43 [393] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3605]    = ( l_43 [394] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3606]    = ( l_43 [395] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3607]    = ( l_43 [396] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3608]    = ( l_43 [397] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3609]    = ( l_43 [398] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[3610]    = ( l_43 [391] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3611]    = ( l_43 [392] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3612]    = ( l_43 [393] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3613]    = ( l_43 [394] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3614]    = ( l_43 [395] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3615]    = ( l_43 [396] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3616]    = ( l_43 [397] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3617]    = ( l_43 [398] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[3618]    = ( l_43 [391] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3619]    = ( l_43 [392] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3620]    = ( l_43 [393] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3621]    = ( l_43 [394] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3622]    = ( l_43 [395] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3623]    = ( l_43 [396] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3624]    = ( l_43 [397] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3625]    = ( l_43 [398] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[3626]    = ( l_43 [391] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3627]    = ( l_43 [392] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3628]    = ( l_43 [393] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3629]    = ( l_43 [394] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3630]    = ( l_43 [395] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3631]    = ( l_43 [396] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3632]    = ( l_43 [397] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3633]    = ( l_43 [398] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[3634]    = ( l_43 [391] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3635]    = ( l_43 [392] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3636]    = ( l_43 [393] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3637]    = ( l_43 [394] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3638]    = ( l_43 [395] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3639]    = ( l_43 [396] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3640]    = ( l_43 [397] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3641]    = ( l_43 [398] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[3642]    = ( l_43 [391] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3643]    = ( l_43 [392] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3644]    = ( l_43 [393] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3645]    = ( l_43 [394] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3646]    = ( l_43 [395] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3647]    = ( l_43 [396] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3648]    = ( l_43 [397] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3649]    = ( l_43 [398] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[3650]    = ( l_43 [391] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3651]    = ( l_43 [392] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3652]    = ( l_43 [393] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3653]    = ( l_43 [394] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3654]    = ( l_43 [395] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3655]    = ( l_43 [396] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3656]    = ( l_43 [397] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3657]    = ( l_43 [398] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[3658]    = ( l_43 [391] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3659]    = ( l_43 [392] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3660]    = ( l_43 [393] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3661]    = ( l_43 [394] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3662]    = ( l_43 [395] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3663]    = ( l_43 [396] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3664]    = ( l_43 [397] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3665]    = ( l_43 [398] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[3666]    = ( l_43 [391] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3667]    = ( l_43 [392] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3668]    = ( l_43 [393] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3669]    = ( l_43 [394] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3670]    = ( l_43 [395] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3671]    = ( l_43 [396] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3672]    = ( l_43 [397] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3673]    = ( l_43 [398] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[3674]    = ( l_43 [391] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3675]    = ( l_43 [392] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3676]    = ( l_43 [393] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3677]    = ( l_43 [394] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3678]    = ( l_43 [395] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3679]    = ( l_43 [396] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3680]    = ( l_43 [397] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3681]    = ( l_43 [398] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[3682]    = ( l_43 [391] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3683]    = ( l_43 [392] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3684]    = ( l_43 [393] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3685]    = ( l_43 [394] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3686]    = ( l_43 [395] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3687]    = ( l_43 [396] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3688]    = ( l_43 [397] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3689]    = ( l_43 [398] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[3690]    = ( l_43 [391] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3691]    = ( l_43 [392] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3692]    = ( l_43 [393] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3693]    = ( l_43 [394] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3694]    = ( l_43 [395] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3695]    = ( l_43 [396] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3696]    = ( l_43 [397] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3697]    = ( l_43 [398] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[3698]    = ( l_43 [391] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3699]    = ( l_43 [392] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3700]    = ( l_43 [393] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3701]    = ( l_43 [394] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3702]    = ( l_43 [395] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3703]    = ( l_43 [396] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3704]    = ( l_43 [397] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3705]    = ( l_43 [398] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[3706]    = ( l_43 [391] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3707]    = ( l_43 [392] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3708]    = ( l_43 [393] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3709]    = ( l_43 [394] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3710]    = ( l_43 [395] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3711]    = ( l_43 [396] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3712]    = ( l_43 [397] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3713]    = ( l_43 [398] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[3714]    = ( l_43 [391] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3715]    = ( l_43 [392] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3716]    = ( l_43 [393] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3717]    = ( l_43 [394] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3718]    = ( l_43 [395] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3719]    = ( l_43 [396] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3720]    = ( l_43 [397] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3721]    = ( l_43 [398] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[3722]    = ( l_43 [391] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3723]    = ( l_43 [392] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3724]    = ( l_43 [393] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3725]    = ( l_43 [394] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3726]    = ( l_43 [395] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3727]    = ( l_43 [396] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3728]    = ( l_43 [397] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3729]    = ( l_43 [398] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[3730]    = ( l_43 [391] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3731]    = ( l_43 [392] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3732]    = ( l_43 [393] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3733]    = ( l_43 [394] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3734]    = ( l_43 [395] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3735]    = ( l_43 [396] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3736]    = ( l_43 [397] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3737]    = ( l_43 [398] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[3738]    = ( l_43 [391] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3739]    = ( l_43 [392] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3740]    = ( l_43 [393] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3741]    = ( l_43 [394] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3742]    = ( l_43 [395] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3743]    = ( l_43 [396] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3744]    = ( l_43 [397] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3745]    = ( l_43 [398] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[3746]    = ( l_43 [391] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3747]    = ( l_43 [392] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3748]    = ( l_43 [393] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3749]    = ( l_43 [394] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3750]    = ( l_43 [395] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3751]    = ( l_43 [396] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3752]    = ( l_43 [397] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3753]    = ( l_43 [398] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[3754]    = ( l_43 [391] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3755]    = ( l_43 [392] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3756]    = ( l_43 [393] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3757]    = ( l_43 [394] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3758]    = ( l_43 [395] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3759]    = ( l_43 [396] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3760]    = ( l_43 [397] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3761]    = ( l_43 [398] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[3762]    = ( l_43 [391] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3763]    = ( l_43 [392] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3764]    = ( l_43 [393] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3765]    = ( l_43 [394] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3766]    = ( l_43 [395] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3767]    = ( l_43 [396] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3768]    = ( l_43 [397] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3769]    = ( l_43 [398] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[3770]    = ( l_43 [391] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3771]    = ( l_43 [392] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3772]    = ( l_43 [393] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3773]    = ( l_43 [394] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3774]    = ( l_43 [395] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3775]    = ( l_43 [396] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3776]    = ( l_43 [397] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3777]    = ( l_43 [398] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[3778]    = ( l_43 [391] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3779]    = ( l_43 [392] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3780]    = ( l_43 [393] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3781]    = ( l_43 [394] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3782]    = ( l_43 [395] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3783]    = ( l_43 [396] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3784]    = ( l_43 [397] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3785]    = ( l_43 [398] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[3786]    = ( l_43 [391] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3787]    = ( l_43 [392] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3788]    = ( l_43 [393] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3789]    = ( l_43 [394] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3790]    = ( l_43 [395] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3791]    = ( l_43 [396] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3792]    = ( l_43 [397] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3793]    = ( l_43 [398] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[3794]    = ( l_43 [391] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3795]    = ( l_43 [392] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3796]    = ( l_43 [393] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3797]    = ( l_43 [394] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3798]    = ( l_43 [395] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3799]    = ( l_43 [396] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3800]    = ( l_43 [397] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3801]    = ( l_43 [398] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[3802]    = ( l_43 [391] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3803]    = ( l_43 [392] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3804]    = ( l_43 [393] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3805]    = ( l_43 [394] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3806]    = ( l_43 [395] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3807]    = ( l_43 [396] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3808]    = ( l_43 [397] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3809]    = ( l_43 [398] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[3810]    = ( l_43 [391] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3811]    = ( l_43 [392] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3812]    = ( l_43 [393] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3813]    = ( l_43 [394] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3814]    = ( l_43 [395] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3815]    = ( l_43 [396] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3816]    = ( l_43 [397] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3817]    = ( l_43 [398] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[3818]    = ( l_43 [391] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3819]    = ( l_43 [392] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3820]    = ( l_43 [393] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3821]    = ( l_43 [394] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3822]    = ( l_43 [395] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3823]    = ( l_43 [396] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3824]    = ( l_43 [397] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3825]    = ( l_43 [398] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[3826]    = ( l_43 [391] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3827]    = ( l_43 [392] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3828]    = ( l_43 [393] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3829]    = ( l_43 [394] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3830]    = ( l_43 [395] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3831]    = ( l_43 [396] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3832]    = ( l_43 [397] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3833]    = ( l_43 [398] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[3834]    = ( l_43 [391] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3835]    = ( l_43 [392] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3836]    = ( l_43 [393] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3837]    = ( l_43 [394] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3838]    = ( l_43 [395] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3839]    = ( l_43 [396] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3840]    = ( l_43 [397] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3841]    = ( l_43 [398] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[3842]    = ( l_43 [391] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3843]    = ( l_43 [392] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3844]    = ( l_43 [393] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3845]    = ( l_43 [394] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3846]    = ( l_43 [395] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3847]    = ( l_43 [396] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3848]    = ( l_43 [397] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3849]    = ( l_43 [398] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[3850]    = ( l_43 [391] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3851]    = ( l_43 [392] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3852]    = ( l_43 [393] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3853]    = ( l_43 [394] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3854]    = ( l_43 [395] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3855]    = ( l_43 [396] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3856]    = ( l_43 [397] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3857]    = ( l_43 [398] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[3858]    = ( l_43 [391] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3859]    = ( l_43 [392] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3860]    = ( l_43 [393] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3861]    = ( l_43 [394] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3862]    = ( l_43 [395] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3863]    = ( l_43 [396] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3864]    = ( l_43 [397] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3865]    = ( l_43 [398] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[3866]    = ( l_43 [391] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3867]    = ( l_43 [392] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3868]    = ( l_43 [393] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3869]    = ( l_43 [394] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3870]    = ( l_43 [395] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3871]    = ( l_43 [396] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3872]    = ( l_43 [397] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3873]    = ( l_43 [398] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[3874]    = ( l_43 [391] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3875]    = ( l_43 [392] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3876]    = ( l_43 [393] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3877]    = ( l_43 [394] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3878]    = ( l_43 [395] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3879]    = ( l_43 [396] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3880]    = ( l_43 [397] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3881]    = ( l_43 [398] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[3882]    = ( l_43 [391] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3883]    = ( l_43 [392] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3884]    = ( l_43 [393] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3885]    = ( l_43 [394] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3886]    = ( l_43 [395] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3887]    = ( l_43 [396] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3888]    = ( l_43 [397] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3889]    = ( l_43 [398] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[3890]    = ( l_43 [391] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3891]    = ( l_43 [392] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3892]    = ( l_43 [393] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3893]    = ( l_43 [394] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3894]    = ( l_43 [395] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3895]    = ( l_43 [396] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3896]    = ( l_43 [397] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3897]    = ( l_43 [398] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[3898]    = ( l_43 [391] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3899]    = ( l_43 [392] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3900]    = ( l_43 [393] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3901]    = ( l_43 [394] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3902]    = ( l_43 [395] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3903]    = ( l_43 [396] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3904]    = ( l_43 [397] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3905]    = ( l_43 [398] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[3906]    = ( l_43 [391] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3907]    = ( l_43 [392] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3908]    = ( l_43 [393] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3909]    = ( l_43 [394] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3910]    = ( l_43 [395] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3911]    = ( l_43 [396] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3912]    = ( l_43 [397] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3913]    = ( l_43 [398] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[3914]    = ( l_43 [391] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3915]    = ( l_43 [392] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3916]    = ( l_43 [393] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3917]    = ( l_43 [394] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3918]    = ( l_43 [395] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3919]    = ( l_43 [396] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3920]    = ( l_43 [397] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3921]    = ( l_43 [398] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[3922]    = ( l_43 [391] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3923]    = ( l_43 [392] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3924]    = ( l_43 [393] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3925]    = ( l_43 [394] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3926]    = ( l_43 [395] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3927]    = ( l_43 [396] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3928]    = ( l_43 [397] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3929]    = ( l_43 [398] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[3930]    = ( l_43 [391] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3931]    = ( l_43 [392] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3932]    = ( l_43 [393] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3933]    = ( l_43 [394] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3934]    = ( l_43 [395] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3935]    = ( l_43 [396] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3936]    = ( l_43 [397] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3937]    = ( l_43 [398] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[3938]    = ( l_43 [391] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3939]    = ( l_43 [392] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3940]    = ( l_43 [393] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3941]    = ( l_43 [394] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3942]    = ( l_43 [395] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3943]    = ( l_43 [396] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3944]    = ( l_43 [397] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3945]    = ( l_43 [398] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[3946]    = ( l_43 [391] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3947]    = ( l_43 [392] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3948]    = ( l_43 [393] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3949]    = ( l_43 [394] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3950]    = ( l_43 [395] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3951]    = ( l_43 [396] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3952]    = ( l_43 [397] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3953]    = ( l_43 [398] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[3954]    = ( l_43 [391] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3955]    = ( l_43 [392] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3956]    = ( l_43 [393] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3957]    = ( l_43 [394] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3958]    = ( l_43 [395] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3959]    = ( l_43 [396] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3960]    = ( l_43 [397] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3961]    = ( l_43 [398] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[3962]    = ( l_43 [391] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3963]    = ( l_43 [392] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3964]    = ( l_43 [393] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3965]    = ( l_43 [394] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3966]    = ( l_43 [395] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3967]    = ( l_43 [396] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3968]    = ( l_43 [397] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3969]    = ( l_43 [398] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[3970]    = ( l_43 [391] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3971]    = ( l_43 [392] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3972]    = ( l_43 [393] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3973]    = ( l_43 [394] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3974]    = ( l_43 [395] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3975]    = ( l_43 [396] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3976]    = ( l_43 [397] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3977]    = ( l_43 [398] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[3978]    = ( l_43 [391] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3979]    = ( l_43 [392] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3980]    = ( l_43 [393] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3981]    = ( l_43 [394] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3982]    = ( l_43 [395] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3983]    = ( l_43 [396] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3984]    = ( l_43 [397] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3985]    = ( l_43 [398] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[3986]    = ( l_43 [391] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3987]    = ( l_43 [392] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3988]    = ( l_43 [393] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3989]    = ( l_43 [394] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3990]    = ( l_43 [395] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3991]    = ( l_43 [396] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3992]    = ( l_43 [397] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3993]    = ( l_43 [398] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[3994]    = ( l_43 [391] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[3995]    = ( l_43 [392] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[3996]    = ( l_43 [393] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[3997]    = ( l_43 [394] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[3998]    = ( l_43 [395] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[3999]    = ( l_43 [396] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[4000]    = ( l_43 [397] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[4001]    = ( l_43 [398] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[4002]    = ( l_43 [391] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4003]    = ( l_43 [392] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4004]    = ( l_43 [393] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4005]    = ( l_43 [394] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4006]    = ( l_43 [395] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4007]    = ( l_43 [396] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4008]    = ( l_43 [397] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4009]    = ( l_43 [398] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[4010]    = ( l_43 [391] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4011]    = ( l_43 [392] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4012]    = ( l_43 [393] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4013]    = ( l_43 [394] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4014]    = ( l_43 [395] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4015]    = ( l_43 [396] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4016]    = ( l_43 [397] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4017]    = ( l_43 [398] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[4018]    = ( l_43 [391] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4019]    = ( l_43 [392] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4020]    = ( l_43 [393] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4021]    = ( l_43 [394] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4022]    = ( l_43 [395] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4023]    = ( l_43 [396] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4024]    = ( l_43 [397] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4025]    = ( l_43 [398] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[4026]    = ( l_43 [391] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4027]    = ( l_43 [392] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4028]    = ( l_43 [393] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4029]    = ( l_43 [394] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4030]    = ( l_43 [395] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4031]    = ( l_43 [396] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4032]    = ( l_43 [397] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4033]    = ( l_43 [398] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[4034]    = ( l_43 [391] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4035]    = ( l_43 [392] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4036]    = ( l_43 [393] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4037]    = ( l_43 [394] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4038]    = ( l_43 [395] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4039]    = ( l_43 [396] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4040]    = ( l_43 [397] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4041]    = ( l_43 [398] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[4042]    = ( l_43 [391] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4043]    = ( l_43 [392] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4044]    = ( l_43 [393] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4045]    = ( l_43 [394] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4046]    = ( l_43 [395] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4047]    = ( l_43 [396] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4048]    = ( l_43 [397] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4049]    = ( l_43 [398] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[4050]    = ( l_43 [391] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4051]    = ( l_43 [392] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4052]    = ( l_43 [393] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4053]    = ( l_43 [394] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4054]    = ( l_43 [395] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4055]    = ( l_43 [396] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4056]    = ( l_43 [397] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4057]    = ( l_43 [398] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[4058]    = ( l_43 [391] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4059]    = ( l_43 [392] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4060]    = ( l_43 [393] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4061]    = ( l_43 [394] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4062]    = ( l_43 [395] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4063]    = ( l_43 [396] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4064]    = ( l_43 [397] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4065]    = ( l_43 [398] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[4066]    = ( l_43 [391] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4067]    = ( l_43 [392] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4068]    = ( l_43 [393] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4069]    = ( l_43 [394] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4070]    = ( l_43 [395] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4071]    = ( l_43 [396] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4072]    = ( l_43 [397] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4073]    = ( l_43 [398] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[4074]    = ( l_43 [391] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4075]    = ( l_43 [392] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4076]    = ( l_43 [393] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4077]    = ( l_43 [394] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4078]    = ( l_43 [395] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4079]    = ( l_43 [396] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4080]    = ( l_43 [397] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4081]    = ( l_43 [398] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[4082]    = ( l_43 [391] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4083]    = ( l_43 [392] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4084]    = ( l_43 [393] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4085]    = ( l_43 [394] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4086]    = ( l_43 [395] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4087]    = ( l_43 [396] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4088]    = ( l_43 [397] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4089]    = ( l_43 [398] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[4090]    = ( l_43 [391] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4091]    = ( l_43 [392] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4092]    = ( l_43 [393] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4093]    = ( l_43 [394] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4094]    = ( l_43 [395] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4095]    = ( l_43 [396] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4096]    = ( l_43 [397] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4097]    = ( l_43 [398] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[4098]    = ( l_43 [391] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4099]    = ( l_43 [392] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4100]    = ( l_43 [393] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4101]    = ( l_43 [394] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4102]    = ( l_43 [395] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4103]    = ( l_43 [396] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4104]    = ( l_43 [397] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4105]    = ( l_43 [398] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[4106]    = ( l_43 [391] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4107]    = ( l_43 [392] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4108]    = ( l_43 [393] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4109]    = ( l_43 [394] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4110]    = ( l_43 [395] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4111]    = ( l_43 [396] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4112]    = ( l_43 [397] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4113]    = ( l_43 [398] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[4114]    = ( l_43 [391] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4115]    = ( l_43 [392] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4116]    = ( l_43 [393] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4117]    = ( l_43 [394] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4118]    = ( l_43 [395] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4119]    = ( l_43 [396] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4120]    = ( l_43 [397] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4121]    = ( l_43 [398] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[4122]    = ( l_43 [391] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4123]    = ( l_43 [392] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4124]    = ( l_43 [393] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4125]    = ( l_43 [394] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4126]    = ( l_43 [395] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4127]    = ( l_43 [396] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4128]    = ( l_43 [397] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4129]    = ( l_43 [398] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[4130]    = ( l_43 [391] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4131]    = ( l_43 [392] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4132]    = ( l_43 [393] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4133]    = ( l_43 [394] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4134]    = ( l_43 [395] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4135]    = ( l_43 [396] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4136]    = ( l_43 [397] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4137]    = ( l_43 [398] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[4138]    = ( l_43 [391] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4139]    = ( l_43 [392] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4140]    = ( l_43 [393] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4141]    = ( l_43 [394] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4142]    = ( l_43 [395] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4143]    = ( l_43 [396] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4144]    = ( l_43 [397] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4145]    = ( l_43 [398] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[4146]    = ( l_43 [391] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4147]    = ( l_43 [392] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4148]    = ( l_43 [393] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4149]    = ( l_43 [394] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4150]    = ( l_43 [395] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4151]    = ( l_43 [396] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4152]    = ( l_43 [397] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4153]    = ( l_43 [398] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[4154]    = ( l_43 [391] & !i[1703]) | (      i[1703]);
assign l_42[4155]    = ( l_43 [392] & !i[1703]) | (      i[1703]);
assign l_42[4156]    = ( l_43 [393] & !i[1703]) | (      i[1703]);
assign l_42[4157]    = ( l_43 [394] & !i[1703]) | (      i[1703]);
assign l_42[4158]    = ( l_43 [395] & !i[1703]) | (      i[1703]);
assign l_42[4159]    = ( l_43 [396] & !i[1703]) | (      i[1703]);
assign l_42[4160]    = ( l_43 [397] & !i[1703]) | (      i[1703]);
assign l_42[4161]    = ( l_43 [398] & !i[1703]) | (      i[1703]);
assign l_42[4162]    = ( l_43 [399] & !i[1703]);
assign l_42[4163]    = ( l_43 [400] & !i[1703]);
assign l_42[4164]    = ( l_43 [401] & !i[1703]);
assign l_42[4165]    = ( l_43 [402] & !i[1703]);
assign l_42[4166]    = ( l_43 [399] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4167]    = ( l_43 [400] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4168]    = ( l_43 [401] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4169]    = ( l_43 [402] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4170]    = ( l_43 [399] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4171]    = ( l_43 [400] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4172]    = ( l_43 [401] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4173]    = ( l_43 [402] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4174]    = ( l_43 [399] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4175]    = ( l_43 [400] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4176]    = ( l_43 [401] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4177]    = ( l_43 [402] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4178]    = ( l_43 [403] & !i[1703]);
assign l_42[4179]    = ( l_43 [404] & !i[1703]);
assign l_42[4180]    = ( l_43 [405] & !i[1703]);
assign l_42[4181]    = ( l_43 [406] & !i[1703]);
assign l_42[4182]    = ( l_43 [403] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4183]    = ( l_43 [404] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4184]    = ( l_43 [405] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4185]    = ( l_43 [406] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4186]    = ( l_43 [403] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4187]    = ( l_43 [404] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4188]    = ( l_43 [405] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4189]    = ( l_43 [406] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4190]    = ( l_43 [403] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4191]    = ( l_43 [404] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4192]    = ( l_43 [405] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4193]    = ( l_43 [406] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4194]    = ( l_43 [399] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4195]    = ( l_43 [400] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4196]    = ( l_43 [401] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4197]    = ( l_43 [402] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4198]    = ( l_43 [399] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4199]    = ( l_43 [400] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4200]    = ( l_43 [401] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4201]    = ( l_43 [402] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4202]    = ( l_43 [399] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4203]    = ( l_43 [400] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4204]    = ( l_43 [401] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4205]    = ( l_43 [402] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4206]    = ( l_43 [399] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4207]    = ( l_43 [400] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4208]    = ( l_43 [401] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4209]    = ( l_43 [402] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4210]    = ( l_43 [403] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4211]    = ( l_43 [404] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4212]    = ( l_43 [405] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4213]    = ( l_43 [406] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4214]    = ( l_43 [403] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4215]    = ( l_43 [404] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4216]    = ( l_43 [405] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4217]    = ( l_43 [406] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4218]    = ( l_43 [403] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4219]    = ( l_43 [404] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4220]    = ( l_43 [405] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4221]    = ( l_43 [406] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4222]    = ( l_43 [403] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4223]    = ( l_43 [404] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4224]    = ( l_43 [405] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4225]    = ( l_43 [406] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4226]    = ( l_43 [399] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4227]    = ( l_43 [400] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4228]    = ( l_43 [401] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4229]    = ( l_43 [402] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4230]    = ( l_43 [399] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4231]    = ( l_43 [400] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4232]    = ( l_43 [401] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4233]    = ( l_43 [402] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4234]    = ( l_43 [399] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4235]    = ( l_43 [400] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4236]    = ( l_43 [401] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4237]    = ( l_43 [402] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4238]    = ( l_43 [399] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4239]    = ( l_43 [400] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4240]    = ( l_43 [401] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4241]    = ( l_43 [402] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4242]    = ( l_43 [403] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4243]    = ( l_43 [404] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4244]    = ( l_43 [405] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4245]    = ( l_43 [406] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4246]    = ( l_43 [403] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4247]    = ( l_43 [404] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4248]    = ( l_43 [405] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4249]    = ( l_43 [406] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4250]    = ( l_43 [403] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4251]    = ( l_43 [404] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4252]    = ( l_43 [405] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4253]    = ( l_43 [406] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4254]    = ( l_43 [403] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4255]    = ( l_43 [404] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4256]    = ( l_43 [405] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4257]    = ( l_43 [406] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4258]    = ( l_43 [399] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4259]    = ( l_43 [400] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4260]    = ( l_43 [401] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4261]    = ( l_43 [402] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4262]    = ( l_43 [399] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4263]    = ( l_43 [400] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4264]    = ( l_43 [401] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4265]    = ( l_43 [402] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4266]    = ( l_43 [399] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4267]    = ( l_43 [400] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4268]    = ( l_43 [401] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4269]    = ( l_43 [402] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4270]    = ( l_43 [399] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4271]    = ( l_43 [400] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4272]    = ( l_43 [401] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4273]    = ( l_43 [402] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4274]    = ( l_43 [403] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4275]    = ( l_43 [404] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4276]    = ( l_43 [405] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4277]    = ( l_43 [406] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4278]    = ( l_43 [403] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4279]    = ( l_43 [404] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4280]    = ( l_43 [405] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4281]    = ( l_43 [406] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4282]    = ( l_43 [403] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4283]    = ( l_43 [404] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4284]    = ( l_43 [405] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4285]    = ( l_43 [406] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4286]    = ( l_43 [403] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4287]    = ( l_43 [404] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4288]    = ( l_43 [405] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4289]    = ( l_43 [406] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4290]    = ( l_43 [407] & !i[1703]);
assign l_42[4291]    = ( l_43 [408] & !i[1703]);
assign l_42[4292]    = ( l_43 [409] & !i[1703]);
assign l_42[4293]    = ( l_43 [410] & !i[1703]);
assign l_42[4294]    = ( l_43 [407] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4295]    = ( l_43 [408] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4296]    = ( l_43 [409] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4297]    = ( l_43 [410] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4298]    = ( l_43 [407] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4299]    = ( l_43 [408] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4300]    = ( l_43 [409] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4301]    = ( l_43 [410] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4302]    = ( l_43 [407] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4303]    = ( l_43 [408] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4304]    = ( l_43 [409] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4305]    = ( l_43 [410] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4306]    = ( l_43 [411] & !i[1703]);
assign l_42[4307]    = ( l_43 [412] & !i[1703]);
assign l_42[4308]    = ( l_43 [413] & !i[1703]);
assign l_42[4309]    = ( l_43 [414] & !i[1703]);
assign l_42[4310]    = ( l_43 [411] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4311]    = ( l_43 [412] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4312]    = ( l_43 [413] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4313]    = ( l_43 [414] & !i[1703]) | ( l_43 [168] &  i[1703]);
assign l_42[4314]    = ( l_43 [411] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4315]    = ( l_43 [412] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4316]    = ( l_43 [413] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4317]    = ( l_43 [414] & !i[1703]) | ( l_43 [0] &  i[1703]);
assign l_42[4318]    = ( l_43 [411] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4319]    = ( l_43 [412] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4320]    = ( l_43 [413] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4321]    = ( l_43 [414] & !i[1703]) | ( l_43 [169] &  i[1703]);
assign l_42[4322]    = ( l_43 [407] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4323]    = ( l_43 [408] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4324]    = ( l_43 [409] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4325]    = ( l_43 [410] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4326]    = ( l_43 [407] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4327]    = ( l_43 [408] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4328]    = ( l_43 [409] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4329]    = ( l_43 [410] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4330]    = ( l_43 [407] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4331]    = ( l_43 [408] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4332]    = ( l_43 [409] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4333]    = ( l_43 [410] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4334]    = ( l_43 [407] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4335]    = ( l_43 [408] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4336]    = ( l_43 [409] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4337]    = ( l_43 [410] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4338]    = ( l_43 [411] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4339]    = ( l_43 [412] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4340]    = ( l_43 [413] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4341]    = ( l_43 [414] & !i[1703]) | ( l_43 [152] &  i[1703]);
assign l_42[4342]    = ( l_43 [411] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4343]    = ( l_43 [412] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4344]    = ( l_43 [413] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4345]    = ( l_43 [414] & !i[1703]) | ( l_43 [184] &  i[1703]);
assign l_42[4346]    = ( l_43 [411] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4347]    = ( l_43 [412] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4348]    = ( l_43 [413] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4349]    = ( l_43 [414] & !i[1703]) | ( l_43 [153] &  i[1703]);
assign l_42[4350]    = ( l_43 [411] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4351]    = ( l_43 [412] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4352]    = ( l_43 [413] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4353]    = ( l_43 [414] & !i[1703]) | ( l_43 [185] &  i[1703]);
assign l_42[4354]    = ( l_43 [407] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4355]    = ( l_43 [408] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4356]    = ( l_43 [409] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4357]    = ( l_43 [410] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4358]    = ( l_43 [407] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4359]    = ( l_43 [408] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4360]    = ( l_43 [409] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4361]    = ( l_43 [410] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4362]    = ( l_43 [407] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4363]    = ( l_43 [408] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4364]    = ( l_43 [409] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4365]    = ( l_43 [410] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4366]    = ( l_43 [407] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4367]    = ( l_43 [408] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4368]    = ( l_43 [409] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4369]    = ( l_43 [410] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4370]    = ( l_43 [411] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4371]    = ( l_43 [412] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4372]    = ( l_43 [413] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4373]    = ( l_43 [414] & !i[1703]) | ( l_43 [140] &  i[1703]);
assign l_42[4374]    = ( l_43 [411] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4375]    = ( l_43 [412] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4376]    = ( l_43 [413] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4377]    = ( l_43 [414] & !i[1703]) | ( l_43 [172] &  i[1703]);
assign l_42[4378]    = ( l_43 [411] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4379]    = ( l_43 [412] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4380]    = ( l_43 [413] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4381]    = ( l_43 [414] & !i[1703]) | ( l_43 [141] &  i[1703]);
assign l_42[4382]    = ( l_43 [411] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4383]    = ( l_43 [412] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4384]    = ( l_43 [413] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4385]    = ( l_43 [414] & !i[1703]) | ( l_43 [173] &  i[1703]);
assign l_42[4386]    = ( l_43 [407] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4387]    = ( l_43 [408] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4388]    = ( l_43 [409] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4389]    = ( l_43 [410] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4390]    = ( l_43 [407] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4391]    = ( l_43 [408] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4392]    = ( l_43 [409] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4393]    = ( l_43 [410] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4394]    = ( l_43 [407] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4395]    = ( l_43 [408] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4396]    = ( l_43 [409] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4397]    = ( l_43 [410] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4398]    = ( l_43 [407] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4399]    = ( l_43 [408] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4400]    = ( l_43 [409] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4401]    = ( l_43 [410] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4402]    = ( l_43 [411] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4403]    = ( l_43 [412] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4404]    = ( l_43 [413] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4405]    = ( l_43 [414] & !i[1703]) | ( l_43 [156] &  i[1703]);
assign l_42[4406]    = ( l_43 [411] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4407]    = ( l_43 [412] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4408]    = ( l_43 [413] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4409]    = ( l_43 [414] & !i[1703]) | ( l_43 [188] &  i[1703]);
assign l_42[4410]    = ( l_43 [411] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4411]    = ( l_43 [412] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4412]    = ( l_43 [413] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4413]    = ( l_43 [414] & !i[1703]) | ( l_43 [157] &  i[1703]);
assign l_42[4414]    = ( l_43 [411] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4415]    = ( l_43 [412] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4416]    = ( l_43 [413] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4417]    = ( l_43 [414] & !i[1703]) | ( l_43 [189] &  i[1703]);
assign l_42[4418]    = ( l_43 [399] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4419]    = ( l_43 [400] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4420]    = ( l_43 [401] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4421]    = ( l_43 [402] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4422]    = ( l_43 [399] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4423]    = ( l_43 [400] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4424]    = ( l_43 [401] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4425]    = ( l_43 [402] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4426]    = ( l_43 [399] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4427]    = ( l_43 [400] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4428]    = ( l_43 [401] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4429]    = ( l_43 [402] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4430]    = ( l_43 [399] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4431]    = ( l_43 [400] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4432]    = ( l_43 [401] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4433]    = ( l_43 [402] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4434]    = ( l_43 [403] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4435]    = ( l_43 [404] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4436]    = ( l_43 [405] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4437]    = ( l_43 [406] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4438]    = ( l_43 [403] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4439]    = ( l_43 [404] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4440]    = ( l_43 [405] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4441]    = ( l_43 [406] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4442]    = ( l_43 [403] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4443]    = ( l_43 [404] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4444]    = ( l_43 [405] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4445]    = ( l_43 [406] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4446]    = ( l_43 [403] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4447]    = ( l_43 [404] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4448]    = ( l_43 [405] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4449]    = ( l_43 [406] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4450]    = ( l_43 [399] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4451]    = ( l_43 [400] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4452]    = ( l_43 [401] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4453]    = ( l_43 [402] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4454]    = ( l_43 [399] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4455]    = ( l_43 [400] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4456]    = ( l_43 [401] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4457]    = ( l_43 [402] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4458]    = ( l_43 [399] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4459]    = ( l_43 [400] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4460]    = ( l_43 [401] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4461]    = ( l_43 [402] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4462]    = ( l_43 [399] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4463]    = ( l_43 [400] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4464]    = ( l_43 [401] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4465]    = ( l_43 [402] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4466]    = ( l_43 [403] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4467]    = ( l_43 [404] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4468]    = ( l_43 [405] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4469]    = ( l_43 [406] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4470]    = ( l_43 [403] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4471]    = ( l_43 [404] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4472]    = ( l_43 [405] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4473]    = ( l_43 [406] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4474]    = ( l_43 [403] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4475]    = ( l_43 [404] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4476]    = ( l_43 [405] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4477]    = ( l_43 [406] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4478]    = ( l_43 [403] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4479]    = ( l_43 [404] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4480]    = ( l_43 [405] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4481]    = ( l_43 [406] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4482]    = ( l_43 [399] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4483]    = ( l_43 [400] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4484]    = ( l_43 [401] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4485]    = ( l_43 [402] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4486]    = ( l_43 [399] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4487]    = ( l_43 [400] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4488]    = ( l_43 [401] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4489]    = ( l_43 [402] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4490]    = ( l_43 [399] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4491]    = ( l_43 [400] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4492]    = ( l_43 [401] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4493]    = ( l_43 [402] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4494]    = ( l_43 [399] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4495]    = ( l_43 [400] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4496]    = ( l_43 [401] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4497]    = ( l_43 [402] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4498]    = ( l_43 [403] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4499]    = ( l_43 [404] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4500]    = ( l_43 [405] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4501]    = ( l_43 [406] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4502]    = ( l_43 [403] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4503]    = ( l_43 [404] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4504]    = ( l_43 [405] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4505]    = ( l_43 [406] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4506]    = ( l_43 [403] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4507]    = ( l_43 [404] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4508]    = ( l_43 [405] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4509]    = ( l_43 [406] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4510]    = ( l_43 [403] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4511]    = ( l_43 [404] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4512]    = ( l_43 [405] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4513]    = ( l_43 [406] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4514]    = ( l_43 [399] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4515]    = ( l_43 [400] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4516]    = ( l_43 [401] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4517]    = ( l_43 [402] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4518]    = ( l_43 [399] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4519]    = ( l_43 [400] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4520]    = ( l_43 [401] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4521]    = ( l_43 [402] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4522]    = ( l_43 [399] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4523]    = ( l_43 [400] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4524]    = ( l_43 [401] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4525]    = ( l_43 [402] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4526]    = ( l_43 [399] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4527]    = ( l_43 [400] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4528]    = ( l_43 [401] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4529]    = ( l_43 [402] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4530]    = ( l_43 [403] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4531]    = ( l_43 [404] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4532]    = ( l_43 [405] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4533]    = ( l_43 [406] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4534]    = ( l_43 [403] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4535]    = ( l_43 [404] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4536]    = ( l_43 [405] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4537]    = ( l_43 [406] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4538]    = ( l_43 [403] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4539]    = ( l_43 [404] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4540]    = ( l_43 [405] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4541]    = ( l_43 [406] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4542]    = ( l_43 [403] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4543]    = ( l_43 [404] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4544]    = ( l_43 [405] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4545]    = ( l_43 [406] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4546]    = ( l_43 [407] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4547]    = ( l_43 [408] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4548]    = ( l_43 [409] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4549]    = ( l_43 [410] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4550]    = ( l_43 [407] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4551]    = ( l_43 [408] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4552]    = ( l_43 [409] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4553]    = ( l_43 [410] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4554]    = ( l_43 [407] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4555]    = ( l_43 [408] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4556]    = ( l_43 [409] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4557]    = ( l_43 [410] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4558]    = ( l_43 [407] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4559]    = ( l_43 [408] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4560]    = ( l_43 [409] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4561]    = ( l_43 [410] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4562]    = ( l_43 [411] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4563]    = ( l_43 [412] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4564]    = ( l_43 [413] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4565]    = ( l_43 [414] & !i[1703]) | ( l_43 [138] &  i[1703]);
assign l_42[4566]    = ( l_43 [411] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4567]    = ( l_43 [412] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4568]    = ( l_43 [413] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4569]    = ( l_43 [414] & !i[1703]) | ( l_43 [170] &  i[1703]);
assign l_42[4570]    = ( l_43 [411] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4571]    = ( l_43 [412] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4572]    = ( l_43 [413] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4573]    = ( l_43 [414] & !i[1703]) | ( l_43 [139] &  i[1703]);
assign l_42[4574]    = ( l_43 [411] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4575]    = ( l_43 [412] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4576]    = ( l_43 [413] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4577]    = ( l_43 [414] & !i[1703]) | ( l_43 [171] &  i[1703]);
assign l_42[4578]    = ( l_43 [407] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4579]    = ( l_43 [408] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4580]    = ( l_43 [409] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4581]    = ( l_43 [410] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4582]    = ( l_43 [407] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4583]    = ( l_43 [408] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4584]    = ( l_43 [409] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4585]    = ( l_43 [410] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4586]    = ( l_43 [407] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4587]    = ( l_43 [408] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4588]    = ( l_43 [409] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4589]    = ( l_43 [410] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4590]    = ( l_43 [407] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4591]    = ( l_43 [408] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4592]    = ( l_43 [409] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4593]    = ( l_43 [410] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4594]    = ( l_43 [411] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4595]    = ( l_43 [412] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4596]    = ( l_43 [413] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4597]    = ( l_43 [414] & !i[1703]) | ( l_43 [154] &  i[1703]);
assign l_42[4598]    = ( l_43 [411] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4599]    = ( l_43 [412] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4600]    = ( l_43 [413] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4601]    = ( l_43 [414] & !i[1703]) | ( l_43 [186] &  i[1703]);
assign l_42[4602]    = ( l_43 [411] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4603]    = ( l_43 [412] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4604]    = ( l_43 [413] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4605]    = ( l_43 [414] & !i[1703]) | ( l_43 [155] &  i[1703]);
assign l_42[4606]    = ( l_43 [411] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4607]    = ( l_43 [412] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4608]    = ( l_43 [413] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4609]    = ( l_43 [414] & !i[1703]) | ( l_43 [187] &  i[1703]);
assign l_42[4610]    = ( l_43 [407] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4611]    = ( l_43 [408] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4612]    = ( l_43 [409] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4613]    = ( l_43 [410] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4614]    = ( l_43 [407] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4615]    = ( l_43 [408] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4616]    = ( l_43 [409] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4617]    = ( l_43 [410] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4618]    = ( l_43 [407] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4619]    = ( l_43 [408] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4620]    = ( l_43 [409] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4621]    = ( l_43 [410] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4622]    = ( l_43 [407] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4623]    = ( l_43 [408] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4624]    = ( l_43 [409] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4625]    = ( l_43 [410] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4626]    = ( l_43 [411] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4627]    = ( l_43 [412] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4628]    = ( l_43 [413] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4629]    = ( l_43 [414] & !i[1703]) | ( l_43 [142] &  i[1703]);
assign l_42[4630]    = ( l_43 [411] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4631]    = ( l_43 [412] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4632]    = ( l_43 [413] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4633]    = ( l_43 [414] & !i[1703]) | ( l_43 [174] &  i[1703]);
assign l_42[4634]    = ( l_43 [411] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4635]    = ( l_43 [412] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4636]    = ( l_43 [413] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4637]    = ( l_43 [414] & !i[1703]) | ( l_43 [143] &  i[1703]);
assign l_42[4638]    = ( l_43 [411] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4639]    = ( l_43 [412] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4640]    = ( l_43 [413] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4641]    = ( l_43 [414] & !i[1703]) | ( l_43 [175] &  i[1703]);
assign l_42[4642]    = ( l_43 [407] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4643]    = ( l_43 [408] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4644]    = ( l_43 [409] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4645]    = ( l_43 [410] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4646]    = ( l_43 [407] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4647]    = ( l_43 [408] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4648]    = ( l_43 [409] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4649]    = ( l_43 [410] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4650]    = ( l_43 [407] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4651]    = ( l_43 [408] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4652]    = ( l_43 [409] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4653]    = ( l_43 [410] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4654]    = ( l_43 [407] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4655]    = ( l_43 [408] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4656]    = ( l_43 [409] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4657]    = ( l_43 [410] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4658]    = ( l_43 [411] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4659]    = ( l_43 [412] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4660]    = ( l_43 [413] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4661]    = ( l_43 [414] & !i[1703]) | ( l_43 [158] &  i[1703]);
assign l_42[4662]    = ( l_43 [411] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4663]    = ( l_43 [412] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4664]    = ( l_43 [413] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4665]    = ( l_43 [414] & !i[1703]) | ( l_43 [190] &  i[1703]);
assign l_42[4666]    = ( l_43 [411] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4667]    = ( l_43 [412] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4668]    = ( l_43 [413] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4669]    = ( l_43 [414] & !i[1703]) | ( l_43 [159] &  i[1703]);
assign l_42[4670]    = ( l_43 [411] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4671]    = ( l_43 [412] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4672]    = ( l_43 [413] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4673]    = ( l_43 [414] & !i[1703]) | ( l_43 [191] &  i[1703]);
assign l_42[4674]    = ( l_43 [399] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4675]    = ( l_43 [400] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4676]    = ( l_43 [401] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4677]    = ( l_43 [402] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4678]    = ( l_43 [399] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4679]    = ( l_43 [400] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4680]    = ( l_43 [401] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4681]    = ( l_43 [402] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4682]    = ( l_43 [399] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4683]    = ( l_43 [400] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4684]    = ( l_43 [401] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4685]    = ( l_43 [402] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4686]    = ( l_43 [399] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4687]    = ( l_43 [400] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4688]    = ( l_43 [401] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4689]    = ( l_43 [402] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4690]    = ( l_43 [403] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4691]    = ( l_43 [404] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4692]    = ( l_43 [405] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4693]    = ( l_43 [406] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4694]    = ( l_43 [403] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4695]    = ( l_43 [404] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4696]    = ( l_43 [405] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4697]    = ( l_43 [406] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4698]    = ( l_43 [403] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4699]    = ( l_43 [404] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4700]    = ( l_43 [405] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4701]    = ( l_43 [406] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4702]    = ( l_43 [403] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4703]    = ( l_43 [404] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4704]    = ( l_43 [405] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4705]    = ( l_43 [406] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4706]    = ( l_43 [399] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4707]    = ( l_43 [400] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4708]    = ( l_43 [401] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4709]    = ( l_43 [402] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4710]    = ( l_43 [399] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4711]    = ( l_43 [400] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4712]    = ( l_43 [401] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4713]    = ( l_43 [402] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4714]    = ( l_43 [399] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4715]    = ( l_43 [400] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4716]    = ( l_43 [401] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4717]    = ( l_43 [402] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4718]    = ( l_43 [399] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4719]    = ( l_43 [400] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4720]    = ( l_43 [401] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4721]    = ( l_43 [402] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4722]    = ( l_43 [403] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4723]    = ( l_43 [404] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4724]    = ( l_43 [405] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4725]    = ( l_43 [406] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4726]    = ( l_43 [403] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4727]    = ( l_43 [404] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4728]    = ( l_43 [405] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4729]    = ( l_43 [406] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4730]    = ( l_43 [403] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4731]    = ( l_43 [404] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4732]    = ( l_43 [405] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4733]    = ( l_43 [406] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4734]    = ( l_43 [403] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4735]    = ( l_43 [404] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4736]    = ( l_43 [405] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4737]    = ( l_43 [406] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4738]    = ( l_43 [399] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4739]    = ( l_43 [400] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4740]    = ( l_43 [401] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4741]    = ( l_43 [402] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4742]    = ( l_43 [399] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4743]    = ( l_43 [400] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4744]    = ( l_43 [401] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4745]    = ( l_43 [402] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4746]    = ( l_43 [399] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4747]    = ( l_43 [400] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4748]    = ( l_43 [401] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4749]    = ( l_43 [402] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4750]    = ( l_43 [399] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4751]    = ( l_43 [400] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4752]    = ( l_43 [401] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4753]    = ( l_43 [402] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4754]    = ( l_43 [403] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4755]    = ( l_43 [404] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4756]    = ( l_43 [405] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4757]    = ( l_43 [406] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4758]    = ( l_43 [403] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4759]    = ( l_43 [404] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4760]    = ( l_43 [405] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4761]    = ( l_43 [406] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4762]    = ( l_43 [403] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4763]    = ( l_43 [404] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4764]    = ( l_43 [405] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4765]    = ( l_43 [406] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4766]    = ( l_43 [403] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4767]    = ( l_43 [404] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4768]    = ( l_43 [405] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4769]    = ( l_43 [406] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4770]    = ( l_43 [399] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4771]    = ( l_43 [400] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4772]    = ( l_43 [401] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4773]    = ( l_43 [402] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4774]    = ( l_43 [399] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4775]    = ( l_43 [400] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4776]    = ( l_43 [401] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4777]    = ( l_43 [402] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4778]    = ( l_43 [399] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4779]    = ( l_43 [400] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4780]    = ( l_43 [401] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4781]    = ( l_43 [402] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4782]    = ( l_43 [399] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4783]    = ( l_43 [400] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4784]    = ( l_43 [401] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4785]    = ( l_43 [402] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4786]    = ( l_43 [403] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4787]    = ( l_43 [404] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4788]    = ( l_43 [405] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4789]    = ( l_43 [406] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4790]    = ( l_43 [403] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4791]    = ( l_43 [404] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4792]    = ( l_43 [405] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4793]    = ( l_43 [406] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4794]    = ( l_43 [403] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4795]    = ( l_43 [404] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4796]    = ( l_43 [405] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4797]    = ( l_43 [406] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4798]    = ( l_43 [403] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4799]    = ( l_43 [404] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4800]    = ( l_43 [405] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4801]    = ( l_43 [406] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4802]    = ( l_43 [407] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4803]    = ( l_43 [408] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4804]    = ( l_43 [409] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4805]    = ( l_43 [410] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4806]    = ( l_43 [407] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4807]    = ( l_43 [408] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4808]    = ( l_43 [409] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4809]    = ( l_43 [410] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4810]    = ( l_43 [407] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4811]    = ( l_43 [408] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4812]    = ( l_43 [409] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4813]    = ( l_43 [410] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4814]    = ( l_43 [407] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4815]    = ( l_43 [408] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4816]    = ( l_43 [409] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4817]    = ( l_43 [410] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4818]    = ( l_43 [411] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4819]    = ( l_43 [412] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4820]    = ( l_43 [413] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4821]    = ( l_43 [414] & !i[1703]) | ( l_43 [200] &  i[1703]);
assign l_42[4822]    = ( l_43 [411] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4823]    = ( l_43 [412] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4824]    = ( l_43 [413] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4825]    = ( l_43 [414] & !i[1703]) | ( l_43 [232] &  i[1703]);
assign l_42[4826]    = ( l_43 [411] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4827]    = ( l_43 [412] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4828]    = ( l_43 [413] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4829]    = ( l_43 [414] & !i[1703]) | ( l_43 [201] &  i[1703]);
assign l_42[4830]    = ( l_43 [411] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4831]    = ( l_43 [412] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4832]    = ( l_43 [413] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4833]    = ( l_43 [414] & !i[1703]) | ( l_43 [233] &  i[1703]);
assign l_42[4834]    = ( l_43 [407] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4835]    = ( l_43 [408] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4836]    = ( l_43 [409] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4837]    = ( l_43 [410] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4838]    = ( l_43 [407] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4839]    = ( l_43 [408] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4840]    = ( l_43 [409] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4841]    = ( l_43 [410] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4842]    = ( l_43 [407] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4843]    = ( l_43 [408] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4844]    = ( l_43 [409] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4845]    = ( l_43 [410] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4846]    = ( l_43 [407] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4847]    = ( l_43 [408] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4848]    = ( l_43 [409] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4849]    = ( l_43 [410] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4850]    = ( l_43 [411] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4851]    = ( l_43 [412] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4852]    = ( l_43 [413] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4853]    = ( l_43 [414] & !i[1703]) | ( l_43 [216] &  i[1703]);
assign l_42[4854]    = ( l_43 [411] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4855]    = ( l_43 [412] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4856]    = ( l_43 [413] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4857]    = ( l_43 [414] & !i[1703]) | ( l_43 [248] &  i[1703]);
assign l_42[4858]    = ( l_43 [411] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4859]    = ( l_43 [412] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4860]    = ( l_43 [413] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4861]    = ( l_43 [414] & !i[1703]) | ( l_43 [217] &  i[1703]);
assign l_42[4862]    = ( l_43 [411] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4863]    = ( l_43 [412] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4864]    = ( l_43 [413] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4865]    = ( l_43 [414] & !i[1703]) | ( l_43 [249] &  i[1703]);
assign l_42[4866]    = ( l_43 [407] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4867]    = ( l_43 [408] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4868]    = ( l_43 [409] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4869]    = ( l_43 [410] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4870]    = ( l_43 [407] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4871]    = ( l_43 [408] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4872]    = ( l_43 [409] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4873]    = ( l_43 [410] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4874]    = ( l_43 [407] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4875]    = ( l_43 [408] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4876]    = ( l_43 [409] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4877]    = ( l_43 [410] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4878]    = ( l_43 [407] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4879]    = ( l_43 [408] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4880]    = ( l_43 [409] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4881]    = ( l_43 [410] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4882]    = ( l_43 [411] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4883]    = ( l_43 [412] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4884]    = ( l_43 [413] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4885]    = ( l_43 [414] & !i[1703]) | ( l_43 [204] &  i[1703]);
assign l_42[4886]    = ( l_43 [411] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4887]    = ( l_43 [412] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4888]    = ( l_43 [413] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4889]    = ( l_43 [414] & !i[1703]) | ( l_43 [236] &  i[1703]);
assign l_42[4890]    = ( l_43 [411] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4891]    = ( l_43 [412] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4892]    = ( l_43 [413] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4893]    = ( l_43 [414] & !i[1703]) | ( l_43 [205] &  i[1703]);
assign l_42[4894]    = ( l_43 [411] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4895]    = ( l_43 [412] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4896]    = ( l_43 [413] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4897]    = ( l_43 [414] & !i[1703]) | ( l_43 [237] &  i[1703]);
assign l_42[4898]    = ( l_43 [407] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4899]    = ( l_43 [408] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4900]    = ( l_43 [409] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4901]    = ( l_43 [410] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4902]    = ( l_43 [407] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4903]    = ( l_43 [408] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4904]    = ( l_43 [409] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4905]    = ( l_43 [410] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4906]    = ( l_43 [407] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4907]    = ( l_43 [408] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4908]    = ( l_43 [409] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4909]    = ( l_43 [410] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4910]    = ( l_43 [407] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4911]    = ( l_43 [408] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4912]    = ( l_43 [409] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4913]    = ( l_43 [410] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4914]    = ( l_43 [411] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4915]    = ( l_43 [412] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4916]    = ( l_43 [413] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4917]    = ( l_43 [414] & !i[1703]) | ( l_43 [220] &  i[1703]);
assign l_42[4918]    = ( l_43 [411] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4919]    = ( l_43 [412] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4920]    = ( l_43 [413] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4921]    = ( l_43 [414] & !i[1703]) | ( l_43 [252] &  i[1703]);
assign l_42[4922]    = ( l_43 [411] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4923]    = ( l_43 [412] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4924]    = ( l_43 [413] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4925]    = ( l_43 [414] & !i[1703]) | ( l_43 [221] &  i[1703]);
assign l_42[4926]    = ( l_43 [411] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4927]    = ( l_43 [412] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4928]    = ( l_43 [413] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4929]    = ( l_43 [414] & !i[1703]) | ( l_43 [253] &  i[1703]);
assign l_42[4930]    = ( l_43 [399] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4931]    = ( l_43 [400] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4932]    = ( l_43 [401] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4933]    = ( l_43 [402] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4934]    = ( l_43 [399] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4935]    = ( l_43 [400] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4936]    = ( l_43 [401] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4937]    = ( l_43 [402] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4938]    = ( l_43 [399] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4939]    = ( l_43 [400] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4940]    = ( l_43 [401] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4941]    = ( l_43 [402] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4942]    = ( l_43 [399] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4943]    = ( l_43 [400] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4944]    = ( l_43 [401] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4945]    = ( l_43 [402] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4946]    = ( l_43 [403] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4947]    = ( l_43 [404] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4948]    = ( l_43 [405] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4949]    = ( l_43 [406] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[4950]    = ( l_43 [403] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4951]    = ( l_43 [404] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4952]    = ( l_43 [405] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4953]    = ( l_43 [406] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[4954]    = ( l_43 [403] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4955]    = ( l_43 [404] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4956]    = ( l_43 [405] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4957]    = ( l_43 [406] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[4958]    = ( l_43 [403] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4959]    = ( l_43 [404] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4960]    = ( l_43 [405] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4961]    = ( l_43 [406] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[4962]    = ( l_43 [399] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4963]    = ( l_43 [400] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4964]    = ( l_43 [401] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4965]    = ( l_43 [402] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4966]    = ( l_43 [399] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4967]    = ( l_43 [400] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4968]    = ( l_43 [401] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4969]    = ( l_43 [402] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4970]    = ( l_43 [399] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4971]    = ( l_43 [400] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4972]    = ( l_43 [401] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4973]    = ( l_43 [402] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4974]    = ( l_43 [399] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4975]    = ( l_43 [400] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4976]    = ( l_43 [401] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4977]    = ( l_43 [402] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4978]    = ( l_43 [403] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4979]    = ( l_43 [404] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4980]    = ( l_43 [405] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4981]    = ( l_43 [406] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[4982]    = ( l_43 [403] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4983]    = ( l_43 [404] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4984]    = ( l_43 [405] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4985]    = ( l_43 [406] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[4986]    = ( l_43 [403] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4987]    = ( l_43 [404] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4988]    = ( l_43 [405] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4989]    = ( l_43 [406] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[4990]    = ( l_43 [403] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4991]    = ( l_43 [404] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4992]    = ( l_43 [405] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4993]    = ( l_43 [406] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[4994]    = ( l_43 [399] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[4995]    = ( l_43 [400] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[4996]    = ( l_43 [401] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[4997]    = ( l_43 [402] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[4998]    = ( l_43 [399] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[4999]    = ( l_43 [400] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5000]    = ( l_43 [401] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5001]    = ( l_43 [402] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5002]    = ( l_43 [399] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5003]    = ( l_43 [400] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5004]    = ( l_43 [401] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5005]    = ( l_43 [402] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5006]    = ( l_43 [399] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5007]    = ( l_43 [400] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5008]    = ( l_43 [401] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5009]    = ( l_43 [402] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5010]    = ( l_43 [403] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5011]    = ( l_43 [404] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5012]    = ( l_43 [405] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5013]    = ( l_43 [406] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5014]    = ( l_43 [403] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5015]    = ( l_43 [404] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5016]    = ( l_43 [405] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5017]    = ( l_43 [406] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5018]    = ( l_43 [403] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5019]    = ( l_43 [404] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5020]    = ( l_43 [405] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5021]    = ( l_43 [406] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5022]    = ( l_43 [403] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5023]    = ( l_43 [404] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5024]    = ( l_43 [405] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5025]    = ( l_43 [406] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5026]    = ( l_43 [399] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5027]    = ( l_43 [400] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5028]    = ( l_43 [401] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5029]    = ( l_43 [402] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5030]    = ( l_43 [399] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5031]    = ( l_43 [400] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5032]    = ( l_43 [401] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5033]    = ( l_43 [402] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5034]    = ( l_43 [399] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5035]    = ( l_43 [400] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5036]    = ( l_43 [401] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5037]    = ( l_43 [402] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5038]    = ( l_43 [399] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5039]    = ( l_43 [400] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5040]    = ( l_43 [401] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5041]    = ( l_43 [402] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5042]    = ( l_43 [403] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5043]    = ( l_43 [404] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5044]    = ( l_43 [405] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5045]    = ( l_43 [406] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5046]    = ( l_43 [403] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5047]    = ( l_43 [404] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5048]    = ( l_43 [405] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5049]    = ( l_43 [406] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5050]    = ( l_43 [403] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5051]    = ( l_43 [404] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5052]    = ( l_43 [405] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5053]    = ( l_43 [406] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5054]    = ( l_43 [403] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5055]    = ( l_43 [404] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5056]    = ( l_43 [405] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5057]    = ( l_43 [406] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5058]    = ( l_43 [407] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5059]    = ( l_43 [408] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5060]    = ( l_43 [409] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5061]    = ( l_43 [410] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5062]    = ( l_43 [407] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5063]    = ( l_43 [408] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5064]    = ( l_43 [409] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5065]    = ( l_43 [410] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5066]    = ( l_43 [407] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5067]    = ( l_43 [408] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5068]    = ( l_43 [409] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5069]    = ( l_43 [410] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5070]    = ( l_43 [407] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5071]    = ( l_43 [408] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5072]    = ( l_43 [409] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5073]    = ( l_43 [410] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5074]    = ( l_43 [411] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5075]    = ( l_43 [412] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5076]    = ( l_43 [413] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5077]    = ( l_43 [414] & !i[1703]) | ( l_43 [202] &  i[1703]);
assign l_42[5078]    = ( l_43 [411] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5079]    = ( l_43 [412] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5080]    = ( l_43 [413] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5081]    = ( l_43 [414] & !i[1703]) | ( l_43 [234] &  i[1703]);
assign l_42[5082]    = ( l_43 [411] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5083]    = ( l_43 [412] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5084]    = ( l_43 [413] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5085]    = ( l_43 [414] & !i[1703]) | ( l_43 [203] &  i[1703]);
assign l_42[5086]    = ( l_43 [411] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5087]    = ( l_43 [412] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5088]    = ( l_43 [413] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5089]    = ( l_43 [414] & !i[1703]) | ( l_43 [235] &  i[1703]);
assign l_42[5090]    = ( l_43 [407] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5091]    = ( l_43 [408] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5092]    = ( l_43 [409] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5093]    = ( l_43 [410] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5094]    = ( l_43 [407] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5095]    = ( l_43 [408] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5096]    = ( l_43 [409] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5097]    = ( l_43 [410] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5098]    = ( l_43 [407] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5099]    = ( l_43 [408] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5100]    = ( l_43 [409] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5101]    = ( l_43 [410] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5102]    = ( l_43 [407] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5103]    = ( l_43 [408] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5104]    = ( l_43 [409] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5105]    = ( l_43 [410] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5106]    = ( l_43 [411] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5107]    = ( l_43 [412] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5108]    = ( l_43 [413] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5109]    = ( l_43 [414] & !i[1703]) | ( l_43 [218] &  i[1703]);
assign l_42[5110]    = ( l_43 [411] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5111]    = ( l_43 [412] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5112]    = ( l_43 [413] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5113]    = ( l_43 [414] & !i[1703]) | ( l_43 [250] &  i[1703]);
assign l_42[5114]    = ( l_43 [411] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5115]    = ( l_43 [412] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5116]    = ( l_43 [413] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5117]    = ( l_43 [414] & !i[1703]) | ( l_43 [219] &  i[1703]);
assign l_42[5118]    = ( l_43 [411] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5119]    = ( l_43 [412] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5120]    = ( l_43 [413] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5121]    = ( l_43 [414] & !i[1703]) | ( l_43 [251] &  i[1703]);
assign l_42[5122]    = ( l_43 [407] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5123]    = ( l_43 [408] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5124]    = ( l_43 [409] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5125]    = ( l_43 [410] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5126]    = ( l_43 [407] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5127]    = ( l_43 [408] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5128]    = ( l_43 [409] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5129]    = ( l_43 [410] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5130]    = ( l_43 [407] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5131]    = ( l_43 [408] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5132]    = ( l_43 [409] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5133]    = ( l_43 [410] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5134]    = ( l_43 [407] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5135]    = ( l_43 [408] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5136]    = ( l_43 [409] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5137]    = ( l_43 [410] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5138]    = ( l_43 [411] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5139]    = ( l_43 [412] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5140]    = ( l_43 [413] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5141]    = ( l_43 [414] & !i[1703]) | ( l_43 [206] &  i[1703]);
assign l_42[5142]    = ( l_43 [411] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5143]    = ( l_43 [412] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5144]    = ( l_43 [413] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5145]    = ( l_43 [414] & !i[1703]) | ( l_43 [238] &  i[1703]);
assign l_42[5146]    = ( l_43 [411] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5147]    = ( l_43 [412] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5148]    = ( l_43 [413] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5149]    = ( l_43 [414] & !i[1703]) | ( l_43 [207] &  i[1703]);
assign l_42[5150]    = ( l_43 [411] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5151]    = ( l_43 [412] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5152]    = ( l_43 [413] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5153]    = ( l_43 [414] & !i[1703]) | ( l_43 [239] &  i[1703]);
assign l_42[5154]    = ( l_43 [407] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5155]    = ( l_43 [408] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5156]    = ( l_43 [409] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5157]    = ( l_43 [410] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5158]    = ( l_43 [407] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5159]    = ( l_43 [408] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5160]    = ( l_43 [409] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5161]    = ( l_43 [410] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5162]    = ( l_43 [407] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5163]    = ( l_43 [408] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5164]    = ( l_43 [409] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5165]    = ( l_43 [410] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5166]    = ( l_43 [407] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5167]    = ( l_43 [408] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5168]    = ( l_43 [409] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5169]    = ( l_43 [410] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5170]    = ( l_43 [411] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5171]    = ( l_43 [412] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5172]    = ( l_43 [413] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5173]    = ( l_43 [414] & !i[1703]) | ( l_43 [222] &  i[1703]);
assign l_42[5174]    = ( l_43 [411] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5175]    = ( l_43 [412] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5176]    = ( l_43 [413] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5177]    = ( l_43 [414] & !i[1703]) | ( l_43 [254] &  i[1703]);
assign l_42[5178]    = ( l_43 [411] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5179]    = ( l_43 [412] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5180]    = ( l_43 [413] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5181]    = ( l_43 [414] & !i[1703]) | ( l_43 [223] &  i[1703]);
assign l_42[5182]    = ( l_43 [411] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5183]    = ( l_43 [412] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5184]    = ( l_43 [413] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5185]    = ( l_43 [414] & !i[1703]) | ( l_43 [255] &  i[1703]);
assign l_42[5186]    = ( l_43 [399] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5187]    = ( l_43 [400] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5188]    = ( l_43 [401] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5189]    = ( l_43 [402] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5190]    = ( l_43 [399] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5191]    = ( l_43 [400] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5192]    = ( l_43 [401] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5193]    = ( l_43 [402] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5194]    = ( l_43 [399] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5195]    = ( l_43 [400] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5196]    = ( l_43 [401] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5197]    = ( l_43 [402] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5198]    = ( l_43 [399] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5199]    = ( l_43 [400] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5200]    = ( l_43 [401] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5201]    = ( l_43 [402] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5202]    = ( l_43 [403] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5203]    = ( l_43 [404] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5204]    = ( l_43 [405] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5205]    = ( l_43 [406] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5206]    = ( l_43 [403] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5207]    = ( l_43 [404] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5208]    = ( l_43 [405] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5209]    = ( l_43 [406] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5210]    = ( l_43 [403] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5211]    = ( l_43 [404] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5212]    = ( l_43 [405] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5213]    = ( l_43 [406] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5214]    = ( l_43 [403] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5215]    = ( l_43 [404] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5216]    = ( l_43 [405] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5217]    = ( l_43 [406] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5218]    = ( l_43 [399] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5219]    = ( l_43 [400] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5220]    = ( l_43 [401] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5221]    = ( l_43 [402] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5222]    = ( l_43 [399] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5223]    = ( l_43 [400] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5224]    = ( l_43 [401] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5225]    = ( l_43 [402] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5226]    = ( l_43 [399] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5227]    = ( l_43 [400] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5228]    = ( l_43 [401] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5229]    = ( l_43 [402] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5230]    = ( l_43 [399] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5231]    = ( l_43 [400] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5232]    = ( l_43 [401] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5233]    = ( l_43 [402] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5234]    = ( l_43 [403] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5235]    = ( l_43 [404] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5236]    = ( l_43 [405] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5237]    = ( l_43 [406] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5238]    = ( l_43 [403] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5239]    = ( l_43 [404] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5240]    = ( l_43 [405] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5241]    = ( l_43 [406] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5242]    = ( l_43 [403] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5243]    = ( l_43 [404] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5244]    = ( l_43 [405] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5245]    = ( l_43 [406] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5246]    = ( l_43 [403] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5247]    = ( l_43 [404] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5248]    = ( l_43 [405] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5249]    = ( l_43 [406] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5250]    = ( l_43 [399] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5251]    = ( l_43 [400] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5252]    = ( l_43 [401] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5253]    = ( l_43 [402] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5254]    = ( l_43 [399] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5255]    = ( l_43 [400] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5256]    = ( l_43 [401] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5257]    = ( l_43 [402] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5258]    = ( l_43 [399] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5259]    = ( l_43 [400] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5260]    = ( l_43 [401] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5261]    = ( l_43 [402] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5262]    = ( l_43 [399] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5263]    = ( l_43 [400] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5264]    = ( l_43 [401] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5265]    = ( l_43 [402] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5266]    = ( l_43 [403] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5267]    = ( l_43 [404] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5268]    = ( l_43 [405] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5269]    = ( l_43 [406] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5270]    = ( l_43 [403] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5271]    = ( l_43 [404] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5272]    = ( l_43 [405] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5273]    = ( l_43 [406] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5274]    = ( l_43 [403] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5275]    = ( l_43 [404] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5276]    = ( l_43 [405] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5277]    = ( l_43 [406] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5278]    = ( l_43 [403] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5279]    = ( l_43 [404] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5280]    = ( l_43 [405] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5281]    = ( l_43 [406] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5282]    = ( l_43 [399] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5283]    = ( l_43 [400] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5284]    = ( l_43 [401] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5285]    = ( l_43 [402] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5286]    = ( l_43 [399] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5287]    = ( l_43 [400] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5288]    = ( l_43 [401] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5289]    = ( l_43 [402] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5290]    = ( l_43 [399] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5291]    = ( l_43 [400] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5292]    = ( l_43 [401] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5293]    = ( l_43 [402] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5294]    = ( l_43 [399] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5295]    = ( l_43 [400] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5296]    = ( l_43 [401] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5297]    = ( l_43 [402] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5298]    = ( l_43 [403] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5299]    = ( l_43 [404] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5300]    = ( l_43 [405] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5301]    = ( l_43 [406] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5302]    = ( l_43 [403] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5303]    = ( l_43 [404] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5304]    = ( l_43 [405] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5305]    = ( l_43 [406] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5306]    = ( l_43 [403] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5307]    = ( l_43 [404] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5308]    = ( l_43 [405] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5309]    = ( l_43 [406] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5310]    = ( l_43 [403] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5311]    = ( l_43 [404] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5312]    = ( l_43 [405] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5313]    = ( l_43 [406] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5314]    = ( l_43 [407] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5315]    = ( l_43 [408] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5316]    = ( l_43 [409] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5317]    = ( l_43 [410] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5318]    = ( l_43 [407] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5319]    = ( l_43 [408] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5320]    = ( l_43 [409] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5321]    = ( l_43 [410] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5322]    = ( l_43 [407] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5323]    = ( l_43 [408] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5324]    = ( l_43 [409] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5325]    = ( l_43 [410] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5326]    = ( l_43 [407] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5327]    = ( l_43 [408] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5328]    = ( l_43 [409] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5329]    = ( l_43 [410] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5330]    = ( l_43 [411] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5331]    = ( l_43 [412] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5332]    = ( l_43 [413] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5333]    = ( l_43 [414] & !i[1703]) | ( l_43 [264] &  i[1703]);
assign l_42[5334]    = ( l_43 [411] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5335]    = ( l_43 [412] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5336]    = ( l_43 [413] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5337]    = ( l_43 [414] & !i[1703]) | ( l_43 [296] &  i[1703]);
assign l_42[5338]    = ( l_43 [411] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5339]    = ( l_43 [412] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5340]    = ( l_43 [413] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5341]    = ( l_43 [414] & !i[1703]) | ( l_43 [265] &  i[1703]);
assign l_42[5342]    = ( l_43 [411] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5343]    = ( l_43 [412] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5344]    = ( l_43 [413] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5345]    = ( l_43 [414] & !i[1703]) | ( l_43 [297] &  i[1703]);
assign l_42[5346]    = ( l_43 [407] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5347]    = ( l_43 [408] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5348]    = ( l_43 [409] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5349]    = ( l_43 [410] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5350]    = ( l_43 [407] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5351]    = ( l_43 [408] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5352]    = ( l_43 [409] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5353]    = ( l_43 [410] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5354]    = ( l_43 [407] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5355]    = ( l_43 [408] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5356]    = ( l_43 [409] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5357]    = ( l_43 [410] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5358]    = ( l_43 [407] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5359]    = ( l_43 [408] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5360]    = ( l_43 [409] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5361]    = ( l_43 [410] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5362]    = ( l_43 [411] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5363]    = ( l_43 [412] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5364]    = ( l_43 [413] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5365]    = ( l_43 [414] & !i[1703]) | ( l_43 [280] &  i[1703]);
assign l_42[5366]    = ( l_43 [411] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5367]    = ( l_43 [412] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5368]    = ( l_43 [413] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5369]    = ( l_43 [414] & !i[1703]) | ( l_43 [312] &  i[1703]);
assign l_42[5370]    = ( l_43 [411] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5371]    = ( l_43 [412] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5372]    = ( l_43 [413] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5373]    = ( l_43 [414] & !i[1703]) | ( l_43 [281] &  i[1703]);
assign l_42[5374]    = ( l_43 [411] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5375]    = ( l_43 [412] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5376]    = ( l_43 [413] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5377]    = ( l_43 [414] & !i[1703]) | ( l_43 [313] &  i[1703]);
assign l_42[5378]    = ( l_43 [407] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5379]    = ( l_43 [408] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5380]    = ( l_43 [409] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5381]    = ( l_43 [410] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5382]    = ( l_43 [407] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5383]    = ( l_43 [408] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5384]    = ( l_43 [409] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5385]    = ( l_43 [410] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5386]    = ( l_43 [407] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5387]    = ( l_43 [408] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5388]    = ( l_43 [409] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5389]    = ( l_43 [410] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5390]    = ( l_43 [407] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5391]    = ( l_43 [408] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5392]    = ( l_43 [409] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5393]    = ( l_43 [410] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5394]    = ( l_43 [411] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5395]    = ( l_43 [412] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5396]    = ( l_43 [413] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5397]    = ( l_43 [414] & !i[1703]) | ( l_43 [268] &  i[1703]);
assign l_42[5398]    = ( l_43 [411] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5399]    = ( l_43 [412] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5400]    = ( l_43 [413] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5401]    = ( l_43 [414] & !i[1703]) | ( l_43 [300] &  i[1703]);
assign l_42[5402]    = ( l_43 [411] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5403]    = ( l_43 [412] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5404]    = ( l_43 [413] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5405]    = ( l_43 [414] & !i[1703]) | ( l_43 [269] &  i[1703]);
assign l_42[5406]    = ( l_43 [411] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5407]    = ( l_43 [412] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5408]    = ( l_43 [413] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5409]    = ( l_43 [414] & !i[1703]) | ( l_43 [301] &  i[1703]);
assign l_42[5410]    = ( l_43 [407] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5411]    = ( l_43 [408] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5412]    = ( l_43 [409] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5413]    = ( l_43 [410] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5414]    = ( l_43 [407] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5415]    = ( l_43 [408] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5416]    = ( l_43 [409] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5417]    = ( l_43 [410] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5418]    = ( l_43 [407] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5419]    = ( l_43 [408] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5420]    = ( l_43 [409] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5421]    = ( l_43 [410] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5422]    = ( l_43 [407] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5423]    = ( l_43 [408] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5424]    = ( l_43 [409] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5425]    = ( l_43 [410] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5426]    = ( l_43 [411] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5427]    = ( l_43 [412] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5428]    = ( l_43 [413] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5429]    = ( l_43 [414] & !i[1703]) | ( l_43 [284] &  i[1703]);
assign l_42[5430]    = ( l_43 [411] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5431]    = ( l_43 [412] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5432]    = ( l_43 [413] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5433]    = ( l_43 [414] & !i[1703]) | ( l_43 [316] &  i[1703]);
assign l_42[5434]    = ( l_43 [411] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5435]    = ( l_43 [412] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5436]    = ( l_43 [413] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5437]    = ( l_43 [414] & !i[1703]) | ( l_43 [285] &  i[1703]);
assign l_42[5438]    = ( l_43 [411] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5439]    = ( l_43 [412] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5440]    = ( l_43 [413] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5441]    = ( l_43 [414] & !i[1703]) | ( l_43 [317] &  i[1703]);
assign l_42[5442]    = ( l_43 [399] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5443]    = ( l_43 [400] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5444]    = ( l_43 [401] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5445]    = ( l_43 [402] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5446]    = ( l_43 [399] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5447]    = ( l_43 [400] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5448]    = ( l_43 [401] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5449]    = ( l_43 [402] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5450]    = ( l_43 [399] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5451]    = ( l_43 [400] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5452]    = ( l_43 [401] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5453]    = ( l_43 [402] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5454]    = ( l_43 [399] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5455]    = ( l_43 [400] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5456]    = ( l_43 [401] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5457]    = ( l_43 [402] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5458]    = ( l_43 [403] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5459]    = ( l_43 [404] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5460]    = ( l_43 [405] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5461]    = ( l_43 [406] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5462]    = ( l_43 [403] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5463]    = ( l_43 [404] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5464]    = ( l_43 [405] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5465]    = ( l_43 [406] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5466]    = ( l_43 [403] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5467]    = ( l_43 [404] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5468]    = ( l_43 [405] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5469]    = ( l_43 [406] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5470]    = ( l_43 [403] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5471]    = ( l_43 [404] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5472]    = ( l_43 [405] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5473]    = ( l_43 [406] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5474]    = ( l_43 [399] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5475]    = ( l_43 [400] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5476]    = ( l_43 [401] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5477]    = ( l_43 [402] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5478]    = ( l_43 [399] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5479]    = ( l_43 [400] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5480]    = ( l_43 [401] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5481]    = ( l_43 [402] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5482]    = ( l_43 [399] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5483]    = ( l_43 [400] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5484]    = ( l_43 [401] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5485]    = ( l_43 [402] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5486]    = ( l_43 [399] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5487]    = ( l_43 [400] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5488]    = ( l_43 [401] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5489]    = ( l_43 [402] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5490]    = ( l_43 [403] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5491]    = ( l_43 [404] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5492]    = ( l_43 [405] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5493]    = ( l_43 [406] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5494]    = ( l_43 [403] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5495]    = ( l_43 [404] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5496]    = ( l_43 [405] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5497]    = ( l_43 [406] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5498]    = ( l_43 [403] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5499]    = ( l_43 [404] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5500]    = ( l_43 [405] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5501]    = ( l_43 [406] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5502]    = ( l_43 [403] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5503]    = ( l_43 [404] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5504]    = ( l_43 [405] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5505]    = ( l_43 [406] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5506]    = ( l_43 [399] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5507]    = ( l_43 [400] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5508]    = ( l_43 [401] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5509]    = ( l_43 [402] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5510]    = ( l_43 [399] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5511]    = ( l_43 [400] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5512]    = ( l_43 [401] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5513]    = ( l_43 [402] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5514]    = ( l_43 [399] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5515]    = ( l_43 [400] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5516]    = ( l_43 [401] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5517]    = ( l_43 [402] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5518]    = ( l_43 [399] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5519]    = ( l_43 [400] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5520]    = ( l_43 [401] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5521]    = ( l_43 [402] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5522]    = ( l_43 [403] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5523]    = ( l_43 [404] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5524]    = ( l_43 [405] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5525]    = ( l_43 [406] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5526]    = ( l_43 [403] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5527]    = ( l_43 [404] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5528]    = ( l_43 [405] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5529]    = ( l_43 [406] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5530]    = ( l_43 [403] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5531]    = ( l_43 [404] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5532]    = ( l_43 [405] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5533]    = ( l_43 [406] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5534]    = ( l_43 [403] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5535]    = ( l_43 [404] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5536]    = ( l_43 [405] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5537]    = ( l_43 [406] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5538]    = ( l_43 [399] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5539]    = ( l_43 [400] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5540]    = ( l_43 [401] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5541]    = ( l_43 [402] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5542]    = ( l_43 [399] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5543]    = ( l_43 [400] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5544]    = ( l_43 [401] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5545]    = ( l_43 [402] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5546]    = ( l_43 [399] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5547]    = ( l_43 [400] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5548]    = ( l_43 [401] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5549]    = ( l_43 [402] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5550]    = ( l_43 [399] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5551]    = ( l_43 [400] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5552]    = ( l_43 [401] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5553]    = ( l_43 [402] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5554]    = ( l_43 [403] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5555]    = ( l_43 [404] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5556]    = ( l_43 [405] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5557]    = ( l_43 [406] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5558]    = ( l_43 [403] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5559]    = ( l_43 [404] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5560]    = ( l_43 [405] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5561]    = ( l_43 [406] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5562]    = ( l_43 [403] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5563]    = ( l_43 [404] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5564]    = ( l_43 [405] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5565]    = ( l_43 [406] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5566]    = ( l_43 [403] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5567]    = ( l_43 [404] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5568]    = ( l_43 [405] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5569]    = ( l_43 [406] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5570]    = ( l_43 [407] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5571]    = ( l_43 [408] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5572]    = ( l_43 [409] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5573]    = ( l_43 [410] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5574]    = ( l_43 [407] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5575]    = ( l_43 [408] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5576]    = ( l_43 [409] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5577]    = ( l_43 [410] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5578]    = ( l_43 [407] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5579]    = ( l_43 [408] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5580]    = ( l_43 [409] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5581]    = ( l_43 [410] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5582]    = ( l_43 [407] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5583]    = ( l_43 [408] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5584]    = ( l_43 [409] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5585]    = ( l_43 [410] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5586]    = ( l_43 [411] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5587]    = ( l_43 [412] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5588]    = ( l_43 [413] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5589]    = ( l_43 [414] & !i[1703]) | ( l_43 [266] &  i[1703]);
assign l_42[5590]    = ( l_43 [411] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5591]    = ( l_43 [412] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5592]    = ( l_43 [413] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5593]    = ( l_43 [414] & !i[1703]) | ( l_43 [298] &  i[1703]);
assign l_42[5594]    = ( l_43 [411] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5595]    = ( l_43 [412] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5596]    = ( l_43 [413] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5597]    = ( l_43 [414] & !i[1703]) | ( l_43 [267] &  i[1703]);
assign l_42[5598]    = ( l_43 [411] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5599]    = ( l_43 [412] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5600]    = ( l_43 [413] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5601]    = ( l_43 [414] & !i[1703]) | ( l_43 [299] &  i[1703]);
assign l_42[5602]    = ( l_43 [407] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5603]    = ( l_43 [408] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5604]    = ( l_43 [409] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5605]    = ( l_43 [410] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5606]    = ( l_43 [407] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5607]    = ( l_43 [408] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5608]    = ( l_43 [409] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5609]    = ( l_43 [410] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5610]    = ( l_43 [407] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5611]    = ( l_43 [408] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5612]    = ( l_43 [409] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5613]    = ( l_43 [410] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5614]    = ( l_43 [407] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5615]    = ( l_43 [408] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5616]    = ( l_43 [409] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5617]    = ( l_43 [410] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5618]    = ( l_43 [411] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5619]    = ( l_43 [412] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5620]    = ( l_43 [413] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5621]    = ( l_43 [414] & !i[1703]) | ( l_43 [282] &  i[1703]);
assign l_42[5622]    = ( l_43 [411] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5623]    = ( l_43 [412] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5624]    = ( l_43 [413] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5625]    = ( l_43 [414] & !i[1703]) | ( l_43 [314] &  i[1703]);
assign l_42[5626]    = ( l_43 [411] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5627]    = ( l_43 [412] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5628]    = ( l_43 [413] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5629]    = ( l_43 [414] & !i[1703]) | ( l_43 [283] &  i[1703]);
assign l_42[5630]    = ( l_43 [411] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5631]    = ( l_43 [412] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5632]    = ( l_43 [413] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5633]    = ( l_43 [414] & !i[1703]) | ( l_43 [315] &  i[1703]);
assign l_42[5634]    = ( l_43 [407] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5635]    = ( l_43 [408] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5636]    = ( l_43 [409] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5637]    = ( l_43 [410] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5638]    = ( l_43 [407] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5639]    = ( l_43 [408] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5640]    = ( l_43 [409] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5641]    = ( l_43 [410] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5642]    = ( l_43 [407] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5643]    = ( l_43 [408] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5644]    = ( l_43 [409] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5645]    = ( l_43 [410] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5646]    = ( l_43 [407] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5647]    = ( l_43 [408] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5648]    = ( l_43 [409] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5649]    = ( l_43 [410] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5650]    = ( l_43 [411] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5651]    = ( l_43 [412] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5652]    = ( l_43 [413] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5653]    = ( l_43 [414] & !i[1703]) | ( l_43 [270] &  i[1703]);
assign l_42[5654]    = ( l_43 [411] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5655]    = ( l_43 [412] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5656]    = ( l_43 [413] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5657]    = ( l_43 [414] & !i[1703]) | ( l_43 [302] &  i[1703]);
assign l_42[5658]    = ( l_43 [411] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5659]    = ( l_43 [412] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5660]    = ( l_43 [413] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5661]    = ( l_43 [414] & !i[1703]) | ( l_43 [271] &  i[1703]);
assign l_42[5662]    = ( l_43 [411] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5663]    = ( l_43 [412] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5664]    = ( l_43 [413] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5665]    = ( l_43 [414] & !i[1703]) | ( l_43 [303] &  i[1703]);
assign l_42[5666]    = ( l_43 [407] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5667]    = ( l_43 [408] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5668]    = ( l_43 [409] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5669]    = ( l_43 [410] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5670]    = ( l_43 [407] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5671]    = ( l_43 [408] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5672]    = ( l_43 [409] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5673]    = ( l_43 [410] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5674]    = ( l_43 [407] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5675]    = ( l_43 [408] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5676]    = ( l_43 [409] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5677]    = ( l_43 [410] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5678]    = ( l_43 [407] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5679]    = ( l_43 [408] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5680]    = ( l_43 [409] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5681]    = ( l_43 [410] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5682]    = ( l_43 [411] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5683]    = ( l_43 [412] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5684]    = ( l_43 [413] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5685]    = ( l_43 [414] & !i[1703]) | ( l_43 [286] &  i[1703]);
assign l_42[5686]    = ( l_43 [411] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5687]    = ( l_43 [412] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5688]    = ( l_43 [413] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5689]    = ( l_43 [414] & !i[1703]) | ( l_43 [318] &  i[1703]);
assign l_42[5690]    = ( l_43 [411] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5691]    = ( l_43 [412] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5692]    = ( l_43 [413] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5693]    = ( l_43 [414] & !i[1703]) | ( l_43 [287] &  i[1703]);
assign l_42[5694]    = ( l_43 [411] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5695]    = ( l_43 [412] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5696]    = ( l_43 [413] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5697]    = ( l_43 [414] & !i[1703]) | ( l_43 [319] &  i[1703]);
assign l_42[5698]    = ( l_43 [399] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5699]    = ( l_43 [400] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5700]    = ( l_43 [401] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5701]    = ( l_43 [402] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5702]    = ( l_43 [399] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5703]    = ( l_43 [400] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5704]    = ( l_43 [401] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5705]    = ( l_43 [402] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5706]    = ( l_43 [399] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5707]    = ( l_43 [400] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5708]    = ( l_43 [401] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5709]    = ( l_43 [402] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5710]    = ( l_43 [399] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5711]    = ( l_43 [400] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5712]    = ( l_43 [401] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5713]    = ( l_43 [402] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5714]    = ( l_43 [403] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5715]    = ( l_43 [404] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5716]    = ( l_43 [405] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5717]    = ( l_43 [406] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5718]    = ( l_43 [403] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5719]    = ( l_43 [404] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5720]    = ( l_43 [405] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5721]    = ( l_43 [406] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5722]    = ( l_43 [403] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5723]    = ( l_43 [404] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5724]    = ( l_43 [405] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5725]    = ( l_43 [406] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5726]    = ( l_43 [403] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5727]    = ( l_43 [404] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5728]    = ( l_43 [405] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5729]    = ( l_43 [406] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5730]    = ( l_43 [399] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5731]    = ( l_43 [400] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5732]    = ( l_43 [401] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5733]    = ( l_43 [402] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5734]    = ( l_43 [399] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5735]    = ( l_43 [400] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5736]    = ( l_43 [401] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5737]    = ( l_43 [402] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5738]    = ( l_43 [399] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5739]    = ( l_43 [400] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5740]    = ( l_43 [401] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5741]    = ( l_43 [402] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5742]    = ( l_43 [399] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5743]    = ( l_43 [400] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5744]    = ( l_43 [401] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5745]    = ( l_43 [402] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5746]    = ( l_43 [403] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5747]    = ( l_43 [404] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5748]    = ( l_43 [405] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5749]    = ( l_43 [406] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5750]    = ( l_43 [403] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5751]    = ( l_43 [404] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5752]    = ( l_43 [405] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5753]    = ( l_43 [406] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5754]    = ( l_43 [403] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5755]    = ( l_43 [404] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5756]    = ( l_43 [405] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5757]    = ( l_43 [406] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5758]    = ( l_43 [403] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5759]    = ( l_43 [404] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5760]    = ( l_43 [405] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5761]    = ( l_43 [406] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5762]    = ( l_43 [399] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5763]    = ( l_43 [400] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5764]    = ( l_43 [401] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5765]    = ( l_43 [402] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5766]    = ( l_43 [399] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5767]    = ( l_43 [400] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5768]    = ( l_43 [401] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5769]    = ( l_43 [402] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5770]    = ( l_43 [399] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5771]    = ( l_43 [400] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5772]    = ( l_43 [401] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5773]    = ( l_43 [402] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5774]    = ( l_43 [399] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5775]    = ( l_43 [400] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5776]    = ( l_43 [401] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5777]    = ( l_43 [402] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5778]    = ( l_43 [403] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5779]    = ( l_43 [404] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5780]    = ( l_43 [405] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5781]    = ( l_43 [406] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5782]    = ( l_43 [403] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5783]    = ( l_43 [404] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5784]    = ( l_43 [405] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5785]    = ( l_43 [406] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5786]    = ( l_43 [403] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5787]    = ( l_43 [404] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5788]    = ( l_43 [405] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5789]    = ( l_43 [406] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5790]    = ( l_43 [403] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5791]    = ( l_43 [404] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5792]    = ( l_43 [405] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5793]    = ( l_43 [406] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5794]    = ( l_43 [399] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5795]    = ( l_43 [400] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5796]    = ( l_43 [401] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5797]    = ( l_43 [402] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5798]    = ( l_43 [399] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5799]    = ( l_43 [400] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5800]    = ( l_43 [401] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5801]    = ( l_43 [402] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5802]    = ( l_43 [399] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5803]    = ( l_43 [400] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5804]    = ( l_43 [401] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5805]    = ( l_43 [402] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5806]    = ( l_43 [399] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5807]    = ( l_43 [400] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5808]    = ( l_43 [401] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5809]    = ( l_43 [402] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5810]    = ( l_43 [403] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5811]    = ( l_43 [404] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5812]    = ( l_43 [405] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5813]    = ( l_43 [406] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5814]    = ( l_43 [403] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5815]    = ( l_43 [404] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5816]    = ( l_43 [405] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5817]    = ( l_43 [406] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5818]    = ( l_43 [403] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5819]    = ( l_43 [404] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5820]    = ( l_43 [405] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5821]    = ( l_43 [406] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5822]    = ( l_43 [403] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5823]    = ( l_43 [404] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5824]    = ( l_43 [405] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5825]    = ( l_43 [406] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5826]    = ( l_43 [407] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5827]    = ( l_43 [408] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5828]    = ( l_43 [409] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5829]    = ( l_43 [410] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5830]    = ( l_43 [407] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5831]    = ( l_43 [408] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5832]    = ( l_43 [409] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5833]    = ( l_43 [410] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5834]    = ( l_43 [407] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5835]    = ( l_43 [408] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5836]    = ( l_43 [409] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5837]    = ( l_43 [410] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5838]    = ( l_43 [407] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5839]    = ( l_43 [408] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5840]    = ( l_43 [409] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5841]    = ( l_43 [410] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5842]    = ( l_43 [411] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5843]    = ( l_43 [412] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5844]    = ( l_43 [413] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5845]    = ( l_43 [414] & !i[1703]) | ( l_43 [328] &  i[1703]);
assign l_42[5846]    = ( l_43 [411] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5847]    = ( l_43 [412] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5848]    = ( l_43 [413] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5849]    = ( l_43 [414] & !i[1703]) | ( l_43 [360] &  i[1703]);
assign l_42[5850]    = ( l_43 [411] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5851]    = ( l_43 [412] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5852]    = ( l_43 [413] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5853]    = ( l_43 [414] & !i[1703]) | ( l_43 [329] &  i[1703]);
assign l_42[5854]    = ( l_43 [411] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5855]    = ( l_43 [412] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5856]    = ( l_43 [413] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5857]    = ( l_43 [414] & !i[1703]) | ( l_43 [361] &  i[1703]);
assign l_42[5858]    = ( l_43 [407] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5859]    = ( l_43 [408] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5860]    = ( l_43 [409] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5861]    = ( l_43 [410] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5862]    = ( l_43 [407] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5863]    = ( l_43 [408] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5864]    = ( l_43 [409] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5865]    = ( l_43 [410] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5866]    = ( l_43 [407] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5867]    = ( l_43 [408] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5868]    = ( l_43 [409] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5869]    = ( l_43 [410] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5870]    = ( l_43 [407] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5871]    = ( l_43 [408] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5872]    = ( l_43 [409] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5873]    = ( l_43 [410] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5874]    = ( l_43 [411] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5875]    = ( l_43 [412] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5876]    = ( l_43 [413] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5877]    = ( l_43 [414] & !i[1703]) | ( l_43 [344] &  i[1703]);
assign l_42[5878]    = ( l_43 [411] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5879]    = ( l_43 [412] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5880]    = ( l_43 [413] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5881]    = ( l_43 [414] & !i[1703]) | ( l_43 [376] &  i[1703]);
assign l_42[5882]    = ( l_43 [411] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5883]    = ( l_43 [412] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5884]    = ( l_43 [413] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5885]    = ( l_43 [414] & !i[1703]) | ( l_43 [345] &  i[1703]);
assign l_42[5886]    = ( l_43 [411] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5887]    = ( l_43 [412] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5888]    = ( l_43 [413] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5889]    = ( l_43 [414] & !i[1703]) | ( l_43 [377] &  i[1703]);
assign l_42[5890]    = ( l_43 [407] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5891]    = ( l_43 [408] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5892]    = ( l_43 [409] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5893]    = ( l_43 [410] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5894]    = ( l_43 [407] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5895]    = ( l_43 [408] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5896]    = ( l_43 [409] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5897]    = ( l_43 [410] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5898]    = ( l_43 [407] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5899]    = ( l_43 [408] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5900]    = ( l_43 [409] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5901]    = ( l_43 [410] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5902]    = ( l_43 [407] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5903]    = ( l_43 [408] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5904]    = ( l_43 [409] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5905]    = ( l_43 [410] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5906]    = ( l_43 [411] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5907]    = ( l_43 [412] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5908]    = ( l_43 [413] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5909]    = ( l_43 [414] & !i[1703]) | ( l_43 [332] &  i[1703]);
assign l_42[5910]    = ( l_43 [411] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5911]    = ( l_43 [412] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5912]    = ( l_43 [413] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5913]    = ( l_43 [414] & !i[1703]) | ( l_43 [364] &  i[1703]);
assign l_42[5914]    = ( l_43 [411] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5915]    = ( l_43 [412] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5916]    = ( l_43 [413] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5917]    = ( l_43 [414] & !i[1703]) | ( l_43 [333] &  i[1703]);
assign l_42[5918]    = ( l_43 [411] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5919]    = ( l_43 [412] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5920]    = ( l_43 [413] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5921]    = ( l_43 [414] & !i[1703]) | ( l_43 [365] &  i[1703]);
assign l_42[5922]    = ( l_43 [407] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5923]    = ( l_43 [408] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5924]    = ( l_43 [409] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5925]    = ( l_43 [410] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5926]    = ( l_43 [407] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5927]    = ( l_43 [408] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5928]    = ( l_43 [409] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5929]    = ( l_43 [410] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5930]    = ( l_43 [407] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5931]    = ( l_43 [408] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5932]    = ( l_43 [409] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5933]    = ( l_43 [410] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5934]    = ( l_43 [407] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5935]    = ( l_43 [408] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5936]    = ( l_43 [409] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5937]    = ( l_43 [410] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5938]    = ( l_43 [411] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5939]    = ( l_43 [412] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5940]    = ( l_43 [413] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5941]    = ( l_43 [414] & !i[1703]) | ( l_43 [348] &  i[1703]);
assign l_42[5942]    = ( l_43 [411] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5943]    = ( l_43 [412] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5944]    = ( l_43 [413] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5945]    = ( l_43 [414] & !i[1703]) | ( l_43 [380] &  i[1703]);
assign l_42[5946]    = ( l_43 [411] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5947]    = ( l_43 [412] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5948]    = ( l_43 [413] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5949]    = ( l_43 [414] & !i[1703]) | ( l_43 [349] &  i[1703]);
assign l_42[5950]    = ( l_43 [411] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5951]    = ( l_43 [412] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5952]    = ( l_43 [413] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5953]    = ( l_43 [414] & !i[1703]) | ( l_43 [381] &  i[1703]);
assign l_42[5954]    = ( l_43 [399] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5955]    = ( l_43 [400] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5956]    = ( l_43 [401] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5957]    = ( l_43 [402] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5958]    = ( l_43 [399] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5959]    = ( l_43 [400] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5960]    = ( l_43 [401] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5961]    = ( l_43 [402] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5962]    = ( l_43 [399] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5963]    = ( l_43 [400] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5964]    = ( l_43 [401] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5965]    = ( l_43 [402] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5966]    = ( l_43 [399] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5967]    = ( l_43 [400] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5968]    = ( l_43 [401] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5969]    = ( l_43 [402] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5970]    = ( l_43 [403] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5971]    = ( l_43 [404] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5972]    = ( l_43 [405] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5973]    = ( l_43 [406] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[5974]    = ( l_43 [403] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5975]    = ( l_43 [404] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5976]    = ( l_43 [405] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5977]    = ( l_43 [406] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[5978]    = ( l_43 [403] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5979]    = ( l_43 [404] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5980]    = ( l_43 [405] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5981]    = ( l_43 [406] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[5982]    = ( l_43 [403] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5983]    = ( l_43 [404] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5984]    = ( l_43 [405] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5985]    = ( l_43 [406] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[5986]    = ( l_43 [399] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[5987]    = ( l_43 [400] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[5988]    = ( l_43 [401] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[5989]    = ( l_43 [402] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[5990]    = ( l_43 [399] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[5991]    = ( l_43 [400] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[5992]    = ( l_43 [401] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[5993]    = ( l_43 [402] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[5994]    = ( l_43 [399] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[5995]    = ( l_43 [400] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[5996]    = ( l_43 [401] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[5997]    = ( l_43 [402] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[5998]    = ( l_43 [399] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[5999]    = ( l_43 [400] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6000]    = ( l_43 [401] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6001]    = ( l_43 [402] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6002]    = ( l_43 [403] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6003]    = ( l_43 [404] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6004]    = ( l_43 [405] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6005]    = ( l_43 [406] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6006]    = ( l_43 [403] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6007]    = ( l_43 [404] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6008]    = ( l_43 [405] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6009]    = ( l_43 [406] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6010]    = ( l_43 [403] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6011]    = ( l_43 [404] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6012]    = ( l_43 [405] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6013]    = ( l_43 [406] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6014]    = ( l_43 [403] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6015]    = ( l_43 [404] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6016]    = ( l_43 [405] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6017]    = ( l_43 [406] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6018]    = ( l_43 [399] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6019]    = ( l_43 [400] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6020]    = ( l_43 [401] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6021]    = ( l_43 [402] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6022]    = ( l_43 [399] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6023]    = ( l_43 [400] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6024]    = ( l_43 [401] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6025]    = ( l_43 [402] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6026]    = ( l_43 [399] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6027]    = ( l_43 [400] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6028]    = ( l_43 [401] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6029]    = ( l_43 [402] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6030]    = ( l_43 [399] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6031]    = ( l_43 [400] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6032]    = ( l_43 [401] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6033]    = ( l_43 [402] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6034]    = ( l_43 [403] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6035]    = ( l_43 [404] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6036]    = ( l_43 [405] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6037]    = ( l_43 [406] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6038]    = ( l_43 [403] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6039]    = ( l_43 [404] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6040]    = ( l_43 [405] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6041]    = ( l_43 [406] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6042]    = ( l_43 [403] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6043]    = ( l_43 [404] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6044]    = ( l_43 [405] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6045]    = ( l_43 [406] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6046]    = ( l_43 [403] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6047]    = ( l_43 [404] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6048]    = ( l_43 [405] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6049]    = ( l_43 [406] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6050]    = ( l_43 [399] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6051]    = ( l_43 [400] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6052]    = ( l_43 [401] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6053]    = ( l_43 [402] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6054]    = ( l_43 [399] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6055]    = ( l_43 [400] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6056]    = ( l_43 [401] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6057]    = ( l_43 [402] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6058]    = ( l_43 [399] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6059]    = ( l_43 [400] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6060]    = ( l_43 [401] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6061]    = ( l_43 [402] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6062]    = ( l_43 [399] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6063]    = ( l_43 [400] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6064]    = ( l_43 [401] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6065]    = ( l_43 [402] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6066]    = ( l_43 [403] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6067]    = ( l_43 [404] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6068]    = ( l_43 [405] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6069]    = ( l_43 [406] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6070]    = ( l_43 [403] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6071]    = ( l_43 [404] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6072]    = ( l_43 [405] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6073]    = ( l_43 [406] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6074]    = ( l_43 [403] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6075]    = ( l_43 [404] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6076]    = ( l_43 [405] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6077]    = ( l_43 [406] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6078]    = ( l_43 [403] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6079]    = ( l_43 [404] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6080]    = ( l_43 [405] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6081]    = ( l_43 [406] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6082]    = ( l_43 [407] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6083]    = ( l_43 [408] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6084]    = ( l_43 [409] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6085]    = ( l_43 [410] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6086]    = ( l_43 [407] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6087]    = ( l_43 [408] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6088]    = ( l_43 [409] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6089]    = ( l_43 [410] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6090]    = ( l_43 [407] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6091]    = ( l_43 [408] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6092]    = ( l_43 [409] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6093]    = ( l_43 [410] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6094]    = ( l_43 [407] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6095]    = ( l_43 [408] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6096]    = ( l_43 [409] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6097]    = ( l_43 [410] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6098]    = ( l_43 [411] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6099]    = ( l_43 [412] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6100]    = ( l_43 [413] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6101]    = ( l_43 [414] & !i[1703]) | ( l_43 [330] &  i[1703]);
assign l_42[6102]    = ( l_43 [411] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6103]    = ( l_43 [412] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6104]    = ( l_43 [413] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6105]    = ( l_43 [414] & !i[1703]) | ( l_43 [362] &  i[1703]);
assign l_42[6106]    = ( l_43 [411] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6107]    = ( l_43 [412] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6108]    = ( l_43 [413] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6109]    = ( l_43 [414] & !i[1703]) | ( l_43 [331] &  i[1703]);
assign l_42[6110]    = ( l_43 [411] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6111]    = ( l_43 [412] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6112]    = ( l_43 [413] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6113]    = ( l_43 [414] & !i[1703]) | ( l_43 [363] &  i[1703]);
assign l_42[6114]    = ( l_43 [407] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6115]    = ( l_43 [408] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6116]    = ( l_43 [409] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6117]    = ( l_43 [410] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6118]    = ( l_43 [407] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6119]    = ( l_43 [408] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6120]    = ( l_43 [409] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6121]    = ( l_43 [410] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6122]    = ( l_43 [407] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6123]    = ( l_43 [408] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6124]    = ( l_43 [409] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6125]    = ( l_43 [410] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6126]    = ( l_43 [407] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6127]    = ( l_43 [408] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6128]    = ( l_43 [409] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6129]    = ( l_43 [410] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6130]    = ( l_43 [411] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6131]    = ( l_43 [412] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6132]    = ( l_43 [413] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6133]    = ( l_43 [414] & !i[1703]) | ( l_43 [346] &  i[1703]);
assign l_42[6134]    = ( l_43 [411] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6135]    = ( l_43 [412] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6136]    = ( l_43 [413] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6137]    = ( l_43 [414] & !i[1703]) | ( l_43 [378] &  i[1703]);
assign l_42[6138]    = ( l_43 [411] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6139]    = ( l_43 [412] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6140]    = ( l_43 [413] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6141]    = ( l_43 [414] & !i[1703]) | ( l_43 [347] &  i[1703]);
assign l_42[6142]    = ( l_43 [411] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6143]    = ( l_43 [412] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6144]    = ( l_43 [413] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6145]    = ( l_43 [414] & !i[1703]) | ( l_43 [379] &  i[1703]);
assign l_42[6146]    = ( l_43 [407] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6147]    = ( l_43 [408] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6148]    = ( l_43 [409] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6149]    = ( l_43 [410] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6150]    = ( l_43 [407] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6151]    = ( l_43 [408] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6152]    = ( l_43 [409] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6153]    = ( l_43 [410] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6154]    = ( l_43 [407] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6155]    = ( l_43 [408] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6156]    = ( l_43 [409] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6157]    = ( l_43 [410] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6158]    = ( l_43 [407] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6159]    = ( l_43 [408] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6160]    = ( l_43 [409] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6161]    = ( l_43 [410] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6162]    = ( l_43 [411] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6163]    = ( l_43 [412] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6164]    = ( l_43 [413] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6165]    = ( l_43 [414] & !i[1703]) | ( l_43 [334] &  i[1703]);
assign l_42[6166]    = ( l_43 [411] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6167]    = ( l_43 [412] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6168]    = ( l_43 [413] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6169]    = ( l_43 [414] & !i[1703]) | ( l_43 [366] &  i[1703]);
assign l_42[6170]    = ( l_43 [411] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6171]    = ( l_43 [412] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6172]    = ( l_43 [413] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6173]    = ( l_43 [414] & !i[1703]) | ( l_43 [335] &  i[1703]);
assign l_42[6174]    = ( l_43 [411] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6175]    = ( l_43 [412] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6176]    = ( l_43 [413] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6177]    = ( l_43 [414] & !i[1703]) | ( l_43 [367] &  i[1703]);
assign l_42[6178]    = ( l_43 [407] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6179]    = ( l_43 [408] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6180]    = ( l_43 [409] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6181]    = ( l_43 [410] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6182]    = ( l_43 [407] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6183]    = ( l_43 [408] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6184]    = ( l_43 [409] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6185]    = ( l_43 [410] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6186]    = ( l_43 [407] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6187]    = ( l_43 [408] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6188]    = ( l_43 [409] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6189]    = ( l_43 [410] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6190]    = ( l_43 [407] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6191]    = ( l_43 [408] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6192]    = ( l_43 [409] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6193]    = ( l_43 [410] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6194]    = ( l_43 [411] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6195]    = ( l_43 [412] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6196]    = ( l_43 [413] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6197]    = ( l_43 [414] & !i[1703]) | ( l_43 [350] &  i[1703]);
assign l_42[6198]    = ( l_43 [411] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6199]    = ( l_43 [412] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6200]    = ( l_43 [413] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6201]    = ( l_43 [414] & !i[1703]) | ( l_43 [382] &  i[1703]);
assign l_42[6202]    = ( l_43 [411] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6203]    = ( l_43 [412] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6204]    = ( l_43 [413] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6205]    = ( l_43 [414] & !i[1703]) | ( l_43 [351] &  i[1703]);
assign l_42[6206]    = ( l_43 [411] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6207]    = ( l_43 [412] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6208]    = ( l_43 [413] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6209]    = ( l_43 [414] & !i[1703]) | ( l_43 [383] &  i[1703]);
assign l_42[6210]    = ( l_43 [399] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6211]    = ( l_43 [400] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6212]    = ( l_43 [401] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6213]    = ( l_43 [402] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6214]    = ( l_43 [399] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6215]    = ( l_43 [400] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6216]    = ( l_43 [401] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6217]    = ( l_43 [402] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6218]    = ( l_43 [399] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6219]    = ( l_43 [400] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6220]    = ( l_43 [401] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6221]    = ( l_43 [402] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6222]    = ( l_43 [399] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6223]    = ( l_43 [400] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6224]    = ( l_43 [401] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6225]    = ( l_43 [402] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6226]    = ( l_43 [403] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6227]    = ( l_43 [404] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6228]    = ( l_43 [405] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6229]    = ( l_43 [406] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6230]    = ( l_43 [403] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6231]    = ( l_43 [404] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6232]    = ( l_43 [405] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6233]    = ( l_43 [406] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6234]    = ( l_43 [403] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6235]    = ( l_43 [404] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6236]    = ( l_43 [405] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6237]    = ( l_43 [406] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6238]    = ( l_43 [403] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6239]    = ( l_43 [404] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6240]    = ( l_43 [405] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6241]    = ( l_43 [406] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6242]    = ( l_43 [399] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6243]    = ( l_43 [400] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6244]    = ( l_43 [401] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6245]    = ( l_43 [402] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6246]    = ( l_43 [399] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6247]    = ( l_43 [400] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6248]    = ( l_43 [401] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6249]    = ( l_43 [402] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6250]    = ( l_43 [399] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6251]    = ( l_43 [400] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6252]    = ( l_43 [401] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6253]    = ( l_43 [402] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6254]    = ( l_43 [399] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6255]    = ( l_43 [400] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6256]    = ( l_43 [401] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6257]    = ( l_43 [402] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6258]    = ( l_43 [403] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6259]    = ( l_43 [404] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6260]    = ( l_43 [405] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6261]    = ( l_43 [406] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6262]    = ( l_43 [403] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6263]    = ( l_43 [404] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6264]    = ( l_43 [405] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6265]    = ( l_43 [406] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6266]    = ( l_43 [403] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6267]    = ( l_43 [404] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6268]    = ( l_43 [405] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6269]    = ( l_43 [406] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6270]    = ( l_43 [403] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6271]    = ( l_43 [404] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6272]    = ( l_43 [405] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6273]    = ( l_43 [406] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6274]    = ( l_43 [399] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6275]    = ( l_43 [400] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6276]    = ( l_43 [401] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6277]    = ( l_43 [402] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6278]    = ( l_43 [399] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6279]    = ( l_43 [400] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6280]    = ( l_43 [401] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6281]    = ( l_43 [402] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6282]    = ( l_43 [399] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6283]    = ( l_43 [400] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6284]    = ( l_43 [401] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6285]    = ( l_43 [402] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6286]    = ( l_43 [399] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6287]    = ( l_43 [400] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6288]    = ( l_43 [401] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6289]    = ( l_43 [402] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6290]    = ( l_43 [403] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6291]    = ( l_43 [404] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6292]    = ( l_43 [405] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6293]    = ( l_43 [406] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6294]    = ( l_43 [403] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6295]    = ( l_43 [404] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6296]    = ( l_43 [405] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6297]    = ( l_43 [406] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6298]    = ( l_43 [403] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6299]    = ( l_43 [404] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6300]    = ( l_43 [405] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6301]    = ( l_43 [406] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6302]    = ( l_43 [403] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6303]    = ( l_43 [404] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6304]    = ( l_43 [405] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6305]    = ( l_43 [406] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6306]    = ( l_43 [399] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6307]    = ( l_43 [400] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6308]    = ( l_43 [401] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6309]    = ( l_43 [402] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6310]    = ( l_43 [399] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6311]    = ( l_43 [400] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6312]    = ( l_43 [401] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6313]    = ( l_43 [402] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6314]    = ( l_43 [399] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6315]    = ( l_43 [400] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6316]    = ( l_43 [401] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6317]    = ( l_43 [402] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6318]    = ( l_43 [399] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6319]    = ( l_43 [400] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6320]    = ( l_43 [401] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6321]    = ( l_43 [402] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6322]    = ( l_43 [403] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6323]    = ( l_43 [404] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6324]    = ( l_43 [405] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6325]    = ( l_43 [406] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6326]    = ( l_43 [403] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6327]    = ( l_43 [404] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6328]    = ( l_43 [405] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6329]    = ( l_43 [406] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6330]    = ( l_43 [403] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6331]    = ( l_43 [404] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6332]    = ( l_43 [405] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6333]    = ( l_43 [406] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6334]    = ( l_43 [403] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6335]    = ( l_43 [404] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6336]    = ( l_43 [405] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6337]    = ( l_43 [406] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6338]    = ( l_43 [407] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6339]    = ( l_43 [408] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6340]    = ( l_43 [409] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6341]    = ( l_43 [410] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6342]    = ( l_43 [407] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6343]    = ( l_43 [408] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6344]    = ( l_43 [409] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6345]    = ( l_43 [410] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6346]    = ( l_43 [407] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6347]    = ( l_43 [408] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6348]    = ( l_43 [409] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6349]    = ( l_43 [410] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6350]    = ( l_43 [407] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6351]    = ( l_43 [408] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6352]    = ( l_43 [409] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6353]    = ( l_43 [410] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6354]    = ( l_43 [411] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6355]    = ( l_43 [412] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6356]    = ( l_43 [413] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6357]    = ( l_43 [414] & !i[1703]) | ( l_43 [144] &  i[1703]);
assign l_42[6358]    = ( l_43 [411] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6359]    = ( l_43 [412] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6360]    = ( l_43 [413] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6361]    = ( l_43 [414] & !i[1703]) | ( l_43 [176] &  i[1703]);
assign l_42[6362]    = ( l_43 [411] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6363]    = ( l_43 [412] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6364]    = ( l_43 [413] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6365]    = ( l_43 [414] & !i[1703]) | ( l_43 [145] &  i[1703]);
assign l_42[6366]    = ( l_43 [411] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6367]    = ( l_43 [412] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6368]    = ( l_43 [413] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6369]    = ( l_43 [414] & !i[1703]) | ( l_43 [177] &  i[1703]);
assign l_42[6370]    = ( l_43 [407] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6371]    = ( l_43 [408] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6372]    = ( l_43 [409] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6373]    = ( l_43 [410] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6374]    = ( l_43 [407] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6375]    = ( l_43 [408] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6376]    = ( l_43 [409] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6377]    = ( l_43 [410] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6378]    = ( l_43 [407] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6379]    = ( l_43 [408] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6380]    = ( l_43 [409] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6381]    = ( l_43 [410] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6382]    = ( l_43 [407] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6383]    = ( l_43 [408] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6384]    = ( l_43 [409] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6385]    = ( l_43 [410] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6386]    = ( l_43 [411] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6387]    = ( l_43 [412] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6388]    = ( l_43 [413] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6389]    = ( l_43 [414] & !i[1703]) | ( l_43 [160] &  i[1703]);
assign l_42[6390]    = ( l_43 [411] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6391]    = ( l_43 [412] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6392]    = ( l_43 [413] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6393]    = ( l_43 [414] & !i[1703]) | ( l_43 [192] &  i[1703]);
assign l_42[6394]    = ( l_43 [411] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6395]    = ( l_43 [412] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6396]    = ( l_43 [413] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6397]    = ( l_43 [414] & !i[1703]) | ( l_43 [161] &  i[1703]);
assign l_42[6398]    = ( l_43 [411] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6399]    = ( l_43 [412] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6400]    = ( l_43 [413] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6401]    = ( l_43 [414] & !i[1703]) | ( l_43 [193] &  i[1703]);
assign l_42[6402]    = ( l_43 [407] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6403]    = ( l_43 [408] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6404]    = ( l_43 [409] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6405]    = ( l_43 [410] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6406]    = ( l_43 [407] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6407]    = ( l_43 [408] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6408]    = ( l_43 [409] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6409]    = ( l_43 [410] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6410]    = ( l_43 [407] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6411]    = ( l_43 [408] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6412]    = ( l_43 [409] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6413]    = ( l_43 [410] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6414]    = ( l_43 [407] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6415]    = ( l_43 [408] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6416]    = ( l_43 [409] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6417]    = ( l_43 [410] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6418]    = ( l_43 [411] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6419]    = ( l_43 [412] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6420]    = ( l_43 [413] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6421]    = ( l_43 [414] & !i[1703]) | ( l_43 [148] &  i[1703]);
assign l_42[6422]    = ( l_43 [411] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6423]    = ( l_43 [412] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6424]    = ( l_43 [413] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6425]    = ( l_43 [414] & !i[1703]) | ( l_43 [180] &  i[1703]);
assign l_42[6426]    = ( l_43 [411] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6427]    = ( l_43 [412] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6428]    = ( l_43 [413] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6429]    = ( l_43 [414] & !i[1703]) | ( l_43 [149] &  i[1703]);
assign l_42[6430]    = ( l_43 [411] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6431]    = ( l_43 [412] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6432]    = ( l_43 [413] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6433]    = ( l_43 [414] & !i[1703]) | ( l_43 [181] &  i[1703]);
assign l_42[6434]    = ( l_43 [407] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6435]    = ( l_43 [408] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6436]    = ( l_43 [409] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6437]    = ( l_43 [410] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6438]    = ( l_43 [407] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6439]    = ( l_43 [408] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6440]    = ( l_43 [409] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6441]    = ( l_43 [410] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6442]    = ( l_43 [407] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6443]    = ( l_43 [408] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6444]    = ( l_43 [409] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6445]    = ( l_43 [410] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6446]    = ( l_43 [407] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6447]    = ( l_43 [408] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6448]    = ( l_43 [409] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6449]    = ( l_43 [410] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6450]    = ( l_43 [411] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6451]    = ( l_43 [412] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6452]    = ( l_43 [413] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6453]    = ( l_43 [414] & !i[1703]) | ( l_43 [164] &  i[1703]);
assign l_42[6454]    = ( l_43 [411] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6455]    = ( l_43 [412] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6456]    = ( l_43 [413] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6457]    = ( l_43 [414] & !i[1703]) | ( l_43 [196] &  i[1703]);
assign l_42[6458]    = ( l_43 [411] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6459]    = ( l_43 [412] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6460]    = ( l_43 [413] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6461]    = ( l_43 [414] & !i[1703]) | ( l_43 [165] &  i[1703]);
assign l_42[6462]    = ( l_43 [411] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6463]    = ( l_43 [412] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6464]    = ( l_43 [413] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6465]    = ( l_43 [414] & !i[1703]) | ( l_43 [197] &  i[1703]);
assign l_42[6466]    = ( l_43 [399] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6467]    = ( l_43 [400] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6468]    = ( l_43 [401] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6469]    = ( l_43 [402] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6470]    = ( l_43 [399] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6471]    = ( l_43 [400] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6472]    = ( l_43 [401] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6473]    = ( l_43 [402] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6474]    = ( l_43 [399] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6475]    = ( l_43 [400] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6476]    = ( l_43 [401] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6477]    = ( l_43 [402] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6478]    = ( l_43 [399] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6479]    = ( l_43 [400] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6480]    = ( l_43 [401] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6481]    = ( l_43 [402] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6482]    = ( l_43 [403] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6483]    = ( l_43 [404] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6484]    = ( l_43 [405] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6485]    = ( l_43 [406] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6486]    = ( l_43 [403] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6487]    = ( l_43 [404] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6488]    = ( l_43 [405] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6489]    = ( l_43 [406] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6490]    = ( l_43 [403] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6491]    = ( l_43 [404] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6492]    = ( l_43 [405] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6493]    = ( l_43 [406] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6494]    = ( l_43 [403] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6495]    = ( l_43 [404] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6496]    = ( l_43 [405] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6497]    = ( l_43 [406] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6498]    = ( l_43 [399] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6499]    = ( l_43 [400] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6500]    = ( l_43 [401] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6501]    = ( l_43 [402] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6502]    = ( l_43 [399] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6503]    = ( l_43 [400] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6504]    = ( l_43 [401] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6505]    = ( l_43 [402] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6506]    = ( l_43 [399] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6507]    = ( l_43 [400] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6508]    = ( l_43 [401] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6509]    = ( l_43 [402] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6510]    = ( l_43 [399] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6511]    = ( l_43 [400] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6512]    = ( l_43 [401] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6513]    = ( l_43 [402] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6514]    = ( l_43 [403] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6515]    = ( l_43 [404] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6516]    = ( l_43 [405] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6517]    = ( l_43 [406] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6518]    = ( l_43 [403] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6519]    = ( l_43 [404] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6520]    = ( l_43 [405] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6521]    = ( l_43 [406] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6522]    = ( l_43 [403] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6523]    = ( l_43 [404] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6524]    = ( l_43 [405] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6525]    = ( l_43 [406] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6526]    = ( l_43 [403] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6527]    = ( l_43 [404] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6528]    = ( l_43 [405] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6529]    = ( l_43 [406] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6530]    = ( l_43 [399] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6531]    = ( l_43 [400] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6532]    = ( l_43 [401] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6533]    = ( l_43 [402] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6534]    = ( l_43 [399] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6535]    = ( l_43 [400] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6536]    = ( l_43 [401] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6537]    = ( l_43 [402] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6538]    = ( l_43 [399] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6539]    = ( l_43 [400] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6540]    = ( l_43 [401] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6541]    = ( l_43 [402] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6542]    = ( l_43 [399] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6543]    = ( l_43 [400] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6544]    = ( l_43 [401] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6545]    = ( l_43 [402] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6546]    = ( l_43 [403] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6547]    = ( l_43 [404] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6548]    = ( l_43 [405] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6549]    = ( l_43 [406] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6550]    = ( l_43 [403] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6551]    = ( l_43 [404] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6552]    = ( l_43 [405] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6553]    = ( l_43 [406] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6554]    = ( l_43 [403] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6555]    = ( l_43 [404] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6556]    = ( l_43 [405] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6557]    = ( l_43 [406] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6558]    = ( l_43 [403] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6559]    = ( l_43 [404] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6560]    = ( l_43 [405] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6561]    = ( l_43 [406] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6562]    = ( l_43 [399] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6563]    = ( l_43 [400] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6564]    = ( l_43 [401] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6565]    = ( l_43 [402] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6566]    = ( l_43 [399] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6567]    = ( l_43 [400] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6568]    = ( l_43 [401] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6569]    = ( l_43 [402] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6570]    = ( l_43 [399] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6571]    = ( l_43 [400] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6572]    = ( l_43 [401] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6573]    = ( l_43 [402] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6574]    = ( l_43 [399] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6575]    = ( l_43 [400] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6576]    = ( l_43 [401] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6577]    = ( l_43 [402] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6578]    = ( l_43 [403] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6579]    = ( l_43 [404] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6580]    = ( l_43 [405] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6581]    = ( l_43 [406] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6582]    = ( l_43 [403] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6583]    = ( l_43 [404] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6584]    = ( l_43 [405] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6585]    = ( l_43 [406] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6586]    = ( l_43 [403] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6587]    = ( l_43 [404] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6588]    = ( l_43 [405] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6589]    = ( l_43 [406] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6590]    = ( l_43 [403] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6591]    = ( l_43 [404] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6592]    = ( l_43 [405] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6593]    = ( l_43 [406] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6594]    = ( l_43 [407] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6595]    = ( l_43 [408] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6596]    = ( l_43 [409] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6597]    = ( l_43 [410] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6598]    = ( l_43 [407] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6599]    = ( l_43 [408] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6600]    = ( l_43 [409] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6601]    = ( l_43 [410] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6602]    = ( l_43 [407] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6603]    = ( l_43 [408] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6604]    = ( l_43 [409] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6605]    = ( l_43 [410] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6606]    = ( l_43 [407] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6607]    = ( l_43 [408] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6608]    = ( l_43 [409] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6609]    = ( l_43 [410] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6610]    = ( l_43 [411] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6611]    = ( l_43 [412] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6612]    = ( l_43 [413] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6613]    = ( l_43 [414] & !i[1703]) | ( l_43 [146] &  i[1703]);
assign l_42[6614]    = ( l_43 [411] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6615]    = ( l_43 [412] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6616]    = ( l_43 [413] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6617]    = ( l_43 [414] & !i[1703]) | ( l_43 [178] &  i[1703]);
assign l_42[6618]    = ( l_43 [411] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6619]    = ( l_43 [412] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6620]    = ( l_43 [413] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6621]    = ( l_43 [414] & !i[1703]) | ( l_43 [147] &  i[1703]);
assign l_42[6622]    = ( l_43 [411] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6623]    = ( l_43 [412] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6624]    = ( l_43 [413] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6625]    = ( l_43 [414] & !i[1703]) | ( l_43 [179] &  i[1703]);
assign l_42[6626]    = ( l_43 [407] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6627]    = ( l_43 [408] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6628]    = ( l_43 [409] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6629]    = ( l_43 [410] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6630]    = ( l_43 [407] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6631]    = ( l_43 [408] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6632]    = ( l_43 [409] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6633]    = ( l_43 [410] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6634]    = ( l_43 [407] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6635]    = ( l_43 [408] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6636]    = ( l_43 [409] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6637]    = ( l_43 [410] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6638]    = ( l_43 [407] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6639]    = ( l_43 [408] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6640]    = ( l_43 [409] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6641]    = ( l_43 [410] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6642]    = ( l_43 [411] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6643]    = ( l_43 [412] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6644]    = ( l_43 [413] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6645]    = ( l_43 [414] & !i[1703]) | ( l_43 [162] &  i[1703]);
assign l_42[6646]    = ( l_43 [411] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6647]    = ( l_43 [412] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6648]    = ( l_43 [413] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6649]    = ( l_43 [414] & !i[1703]) | ( l_43 [194] &  i[1703]);
assign l_42[6650]    = ( l_43 [411] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6651]    = ( l_43 [412] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6652]    = ( l_43 [413] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6653]    = ( l_43 [414] & !i[1703]) | ( l_43 [163] &  i[1703]);
assign l_42[6654]    = ( l_43 [411] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6655]    = ( l_43 [412] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6656]    = ( l_43 [413] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6657]    = ( l_43 [414] & !i[1703]) | ( l_43 [195] &  i[1703]);
assign l_42[6658]    = ( l_43 [407] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6659]    = ( l_43 [408] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6660]    = ( l_43 [409] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6661]    = ( l_43 [410] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6662]    = ( l_43 [407] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6663]    = ( l_43 [408] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6664]    = ( l_43 [409] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6665]    = ( l_43 [410] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6666]    = ( l_43 [407] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6667]    = ( l_43 [408] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6668]    = ( l_43 [409] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6669]    = ( l_43 [410] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6670]    = ( l_43 [407] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6671]    = ( l_43 [408] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6672]    = ( l_43 [409] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6673]    = ( l_43 [410] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6674]    = ( l_43 [411] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6675]    = ( l_43 [412] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6676]    = ( l_43 [413] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6677]    = ( l_43 [414] & !i[1703]) | ( l_43 [150] &  i[1703]);
assign l_42[6678]    = ( l_43 [411] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6679]    = ( l_43 [412] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6680]    = ( l_43 [413] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6681]    = ( l_43 [414] & !i[1703]) | ( l_43 [182] &  i[1703]);
assign l_42[6682]    = ( l_43 [411] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6683]    = ( l_43 [412] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6684]    = ( l_43 [413] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6685]    = ( l_43 [414] & !i[1703]) | ( l_43 [151] &  i[1703]);
assign l_42[6686]    = ( l_43 [411] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6687]    = ( l_43 [412] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6688]    = ( l_43 [413] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6689]    = ( l_43 [414] & !i[1703]) | ( l_43 [183] &  i[1703]);
assign l_42[6690]    = ( l_43 [407] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6691]    = ( l_43 [408] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6692]    = ( l_43 [409] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6693]    = ( l_43 [410] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6694]    = ( l_43 [407] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6695]    = ( l_43 [408] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6696]    = ( l_43 [409] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6697]    = ( l_43 [410] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6698]    = ( l_43 [407] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6699]    = ( l_43 [408] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6700]    = ( l_43 [409] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6701]    = ( l_43 [410] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6702]    = ( l_43 [407] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6703]    = ( l_43 [408] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6704]    = ( l_43 [409] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6705]    = ( l_43 [410] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6706]    = ( l_43 [411] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6707]    = ( l_43 [412] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6708]    = ( l_43 [413] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6709]    = ( l_43 [414] & !i[1703]) | ( l_43 [166] &  i[1703]);
assign l_42[6710]    = ( l_43 [411] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6711]    = ( l_43 [412] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6712]    = ( l_43 [413] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6713]    = ( l_43 [414] & !i[1703]) | ( l_43 [198] &  i[1703]);
assign l_42[6714]    = ( l_43 [411] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6715]    = ( l_43 [412] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6716]    = ( l_43 [413] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6717]    = ( l_43 [414] & !i[1703]) | ( l_43 [167] &  i[1703]);
assign l_42[6718]    = ( l_43 [411] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6719]    = ( l_43 [412] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6720]    = ( l_43 [413] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6721]    = ( l_43 [414] & !i[1703]) | ( l_43 [199] &  i[1703]);
assign l_42[6722]    = ( l_43 [399] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6723]    = ( l_43 [400] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6724]    = ( l_43 [401] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6725]    = ( l_43 [402] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6726]    = ( l_43 [399] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6727]    = ( l_43 [400] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6728]    = ( l_43 [401] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6729]    = ( l_43 [402] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6730]    = ( l_43 [399] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6731]    = ( l_43 [400] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6732]    = ( l_43 [401] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6733]    = ( l_43 [402] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6734]    = ( l_43 [399] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6735]    = ( l_43 [400] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6736]    = ( l_43 [401] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6737]    = ( l_43 [402] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6738]    = ( l_43 [403] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6739]    = ( l_43 [404] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6740]    = ( l_43 [405] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6741]    = ( l_43 [406] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6742]    = ( l_43 [403] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6743]    = ( l_43 [404] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6744]    = ( l_43 [405] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6745]    = ( l_43 [406] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6746]    = ( l_43 [403] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6747]    = ( l_43 [404] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6748]    = ( l_43 [405] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6749]    = ( l_43 [406] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6750]    = ( l_43 [403] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6751]    = ( l_43 [404] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6752]    = ( l_43 [405] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6753]    = ( l_43 [406] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6754]    = ( l_43 [399] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6755]    = ( l_43 [400] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6756]    = ( l_43 [401] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6757]    = ( l_43 [402] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6758]    = ( l_43 [399] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6759]    = ( l_43 [400] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6760]    = ( l_43 [401] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6761]    = ( l_43 [402] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6762]    = ( l_43 [399] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6763]    = ( l_43 [400] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6764]    = ( l_43 [401] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6765]    = ( l_43 [402] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6766]    = ( l_43 [399] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6767]    = ( l_43 [400] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6768]    = ( l_43 [401] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6769]    = ( l_43 [402] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6770]    = ( l_43 [403] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6771]    = ( l_43 [404] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6772]    = ( l_43 [405] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6773]    = ( l_43 [406] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6774]    = ( l_43 [403] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6775]    = ( l_43 [404] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6776]    = ( l_43 [405] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6777]    = ( l_43 [406] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6778]    = ( l_43 [403] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6779]    = ( l_43 [404] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6780]    = ( l_43 [405] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6781]    = ( l_43 [406] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6782]    = ( l_43 [403] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6783]    = ( l_43 [404] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6784]    = ( l_43 [405] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6785]    = ( l_43 [406] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6786]    = ( l_43 [399] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6787]    = ( l_43 [400] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6788]    = ( l_43 [401] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6789]    = ( l_43 [402] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6790]    = ( l_43 [399] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6791]    = ( l_43 [400] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6792]    = ( l_43 [401] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6793]    = ( l_43 [402] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6794]    = ( l_43 [399] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6795]    = ( l_43 [400] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6796]    = ( l_43 [401] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6797]    = ( l_43 [402] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6798]    = ( l_43 [399] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6799]    = ( l_43 [400] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6800]    = ( l_43 [401] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6801]    = ( l_43 [402] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6802]    = ( l_43 [403] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6803]    = ( l_43 [404] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6804]    = ( l_43 [405] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6805]    = ( l_43 [406] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6806]    = ( l_43 [403] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6807]    = ( l_43 [404] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6808]    = ( l_43 [405] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6809]    = ( l_43 [406] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6810]    = ( l_43 [403] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6811]    = ( l_43 [404] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6812]    = ( l_43 [405] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6813]    = ( l_43 [406] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6814]    = ( l_43 [403] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6815]    = ( l_43 [404] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6816]    = ( l_43 [405] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6817]    = ( l_43 [406] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6818]    = ( l_43 [399] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6819]    = ( l_43 [400] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6820]    = ( l_43 [401] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6821]    = ( l_43 [402] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6822]    = ( l_43 [399] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6823]    = ( l_43 [400] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6824]    = ( l_43 [401] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6825]    = ( l_43 [402] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6826]    = ( l_43 [399] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6827]    = ( l_43 [400] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6828]    = ( l_43 [401] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6829]    = ( l_43 [402] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6830]    = ( l_43 [399] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6831]    = ( l_43 [400] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6832]    = ( l_43 [401] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6833]    = ( l_43 [402] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6834]    = ( l_43 [403] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6835]    = ( l_43 [404] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6836]    = ( l_43 [405] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6837]    = ( l_43 [406] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6838]    = ( l_43 [403] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6839]    = ( l_43 [404] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6840]    = ( l_43 [405] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6841]    = ( l_43 [406] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6842]    = ( l_43 [403] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6843]    = ( l_43 [404] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6844]    = ( l_43 [405] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6845]    = ( l_43 [406] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6846]    = ( l_43 [403] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6847]    = ( l_43 [404] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6848]    = ( l_43 [405] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6849]    = ( l_43 [406] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6850]    = ( l_43 [407] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6851]    = ( l_43 [408] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6852]    = ( l_43 [409] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6853]    = ( l_43 [410] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6854]    = ( l_43 [407] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6855]    = ( l_43 [408] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6856]    = ( l_43 [409] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6857]    = ( l_43 [410] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6858]    = ( l_43 [407] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6859]    = ( l_43 [408] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6860]    = ( l_43 [409] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6861]    = ( l_43 [410] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6862]    = ( l_43 [407] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6863]    = ( l_43 [408] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6864]    = ( l_43 [409] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6865]    = ( l_43 [410] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6866]    = ( l_43 [411] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6867]    = ( l_43 [412] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6868]    = ( l_43 [413] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6869]    = ( l_43 [414] & !i[1703]) | ( l_43 [208] &  i[1703]);
assign l_42[6870]    = ( l_43 [411] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6871]    = ( l_43 [412] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6872]    = ( l_43 [413] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6873]    = ( l_43 [414] & !i[1703]) | ( l_43 [240] &  i[1703]);
assign l_42[6874]    = ( l_43 [411] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6875]    = ( l_43 [412] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6876]    = ( l_43 [413] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6877]    = ( l_43 [414] & !i[1703]) | ( l_43 [209] &  i[1703]);
assign l_42[6878]    = ( l_43 [411] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6879]    = ( l_43 [412] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6880]    = ( l_43 [413] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6881]    = ( l_43 [414] & !i[1703]) | ( l_43 [241] &  i[1703]);
assign l_42[6882]    = ( l_43 [407] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6883]    = ( l_43 [408] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6884]    = ( l_43 [409] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6885]    = ( l_43 [410] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6886]    = ( l_43 [407] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6887]    = ( l_43 [408] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6888]    = ( l_43 [409] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6889]    = ( l_43 [410] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6890]    = ( l_43 [407] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6891]    = ( l_43 [408] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6892]    = ( l_43 [409] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6893]    = ( l_43 [410] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6894]    = ( l_43 [407] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6895]    = ( l_43 [408] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6896]    = ( l_43 [409] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6897]    = ( l_43 [410] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6898]    = ( l_43 [411] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6899]    = ( l_43 [412] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6900]    = ( l_43 [413] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6901]    = ( l_43 [414] & !i[1703]) | ( l_43 [224] &  i[1703]);
assign l_42[6902]    = ( l_43 [411] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6903]    = ( l_43 [412] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6904]    = ( l_43 [413] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6905]    = ( l_43 [414] & !i[1703]) | ( l_43 [256] &  i[1703]);
assign l_42[6906]    = ( l_43 [411] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6907]    = ( l_43 [412] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6908]    = ( l_43 [413] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6909]    = ( l_43 [414] & !i[1703]) | ( l_43 [225] &  i[1703]);
assign l_42[6910]    = ( l_43 [411] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6911]    = ( l_43 [412] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6912]    = ( l_43 [413] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6913]    = ( l_43 [414] & !i[1703]) | ( l_43 [257] &  i[1703]);
assign l_42[6914]    = ( l_43 [407] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6915]    = ( l_43 [408] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6916]    = ( l_43 [409] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6917]    = ( l_43 [410] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6918]    = ( l_43 [407] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6919]    = ( l_43 [408] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6920]    = ( l_43 [409] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6921]    = ( l_43 [410] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6922]    = ( l_43 [407] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6923]    = ( l_43 [408] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6924]    = ( l_43 [409] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6925]    = ( l_43 [410] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6926]    = ( l_43 [407] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6927]    = ( l_43 [408] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6928]    = ( l_43 [409] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6929]    = ( l_43 [410] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6930]    = ( l_43 [411] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6931]    = ( l_43 [412] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6932]    = ( l_43 [413] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6933]    = ( l_43 [414] & !i[1703]) | ( l_43 [212] &  i[1703]);
assign l_42[6934]    = ( l_43 [411] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6935]    = ( l_43 [412] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6936]    = ( l_43 [413] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6937]    = ( l_43 [414] & !i[1703]) | ( l_43 [244] &  i[1703]);
assign l_42[6938]    = ( l_43 [411] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6939]    = ( l_43 [412] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6940]    = ( l_43 [413] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6941]    = ( l_43 [414] & !i[1703]) | ( l_43 [213] &  i[1703]);
assign l_42[6942]    = ( l_43 [411] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6943]    = ( l_43 [412] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6944]    = ( l_43 [413] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6945]    = ( l_43 [414] & !i[1703]) | ( l_43 [245] &  i[1703]);
assign l_42[6946]    = ( l_43 [407] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6947]    = ( l_43 [408] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6948]    = ( l_43 [409] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6949]    = ( l_43 [410] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6950]    = ( l_43 [407] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6951]    = ( l_43 [408] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6952]    = ( l_43 [409] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6953]    = ( l_43 [410] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6954]    = ( l_43 [407] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6955]    = ( l_43 [408] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6956]    = ( l_43 [409] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6957]    = ( l_43 [410] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6958]    = ( l_43 [407] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6959]    = ( l_43 [408] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6960]    = ( l_43 [409] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6961]    = ( l_43 [410] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6962]    = ( l_43 [411] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6963]    = ( l_43 [412] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6964]    = ( l_43 [413] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6965]    = ( l_43 [414] & !i[1703]) | ( l_43 [228] &  i[1703]);
assign l_42[6966]    = ( l_43 [411] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6967]    = ( l_43 [412] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6968]    = ( l_43 [413] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6969]    = ( l_43 [414] & !i[1703]) | ( l_43 [260] &  i[1703]);
assign l_42[6970]    = ( l_43 [411] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6971]    = ( l_43 [412] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6972]    = ( l_43 [413] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6973]    = ( l_43 [414] & !i[1703]) | ( l_43 [229] &  i[1703]);
assign l_42[6974]    = ( l_43 [411] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6975]    = ( l_43 [412] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6976]    = ( l_43 [413] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6977]    = ( l_43 [414] & !i[1703]) | ( l_43 [261] &  i[1703]);
assign l_42[6978]    = ( l_43 [399] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6979]    = ( l_43 [400] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6980]    = ( l_43 [401] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6981]    = ( l_43 [402] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6982]    = ( l_43 [399] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[6983]    = ( l_43 [400] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[6984]    = ( l_43 [401] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[6985]    = ( l_43 [402] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[6986]    = ( l_43 [399] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[6987]    = ( l_43 [400] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[6988]    = ( l_43 [401] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[6989]    = ( l_43 [402] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[6990]    = ( l_43 [399] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[6991]    = ( l_43 [400] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[6992]    = ( l_43 [401] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[6993]    = ( l_43 [402] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[6994]    = ( l_43 [403] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6995]    = ( l_43 [404] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6996]    = ( l_43 [405] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6997]    = ( l_43 [406] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[6998]    = ( l_43 [403] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[6999]    = ( l_43 [404] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7000]    = ( l_43 [405] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7001]    = ( l_43 [406] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7002]    = ( l_43 [403] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7003]    = ( l_43 [404] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7004]    = ( l_43 [405] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7005]    = ( l_43 [406] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7006]    = ( l_43 [403] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7007]    = ( l_43 [404] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7008]    = ( l_43 [405] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7009]    = ( l_43 [406] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7010]    = ( l_43 [399] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7011]    = ( l_43 [400] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7012]    = ( l_43 [401] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7013]    = ( l_43 [402] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7014]    = ( l_43 [399] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7015]    = ( l_43 [400] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7016]    = ( l_43 [401] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7017]    = ( l_43 [402] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7018]    = ( l_43 [399] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7019]    = ( l_43 [400] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7020]    = ( l_43 [401] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7021]    = ( l_43 [402] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7022]    = ( l_43 [399] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7023]    = ( l_43 [400] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7024]    = ( l_43 [401] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7025]    = ( l_43 [402] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7026]    = ( l_43 [403] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7027]    = ( l_43 [404] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7028]    = ( l_43 [405] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7029]    = ( l_43 [406] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7030]    = ( l_43 [403] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7031]    = ( l_43 [404] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7032]    = ( l_43 [405] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7033]    = ( l_43 [406] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7034]    = ( l_43 [403] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7035]    = ( l_43 [404] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7036]    = ( l_43 [405] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7037]    = ( l_43 [406] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7038]    = ( l_43 [403] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7039]    = ( l_43 [404] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7040]    = ( l_43 [405] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7041]    = ( l_43 [406] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7042]    = ( l_43 [399] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7043]    = ( l_43 [400] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7044]    = ( l_43 [401] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7045]    = ( l_43 [402] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7046]    = ( l_43 [399] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7047]    = ( l_43 [400] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7048]    = ( l_43 [401] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7049]    = ( l_43 [402] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7050]    = ( l_43 [399] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7051]    = ( l_43 [400] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7052]    = ( l_43 [401] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7053]    = ( l_43 [402] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7054]    = ( l_43 [399] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7055]    = ( l_43 [400] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7056]    = ( l_43 [401] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7057]    = ( l_43 [402] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7058]    = ( l_43 [403] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7059]    = ( l_43 [404] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7060]    = ( l_43 [405] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7061]    = ( l_43 [406] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7062]    = ( l_43 [403] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7063]    = ( l_43 [404] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7064]    = ( l_43 [405] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7065]    = ( l_43 [406] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7066]    = ( l_43 [403] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7067]    = ( l_43 [404] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7068]    = ( l_43 [405] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7069]    = ( l_43 [406] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7070]    = ( l_43 [403] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7071]    = ( l_43 [404] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7072]    = ( l_43 [405] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7073]    = ( l_43 [406] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7074]    = ( l_43 [399] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7075]    = ( l_43 [400] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7076]    = ( l_43 [401] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7077]    = ( l_43 [402] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7078]    = ( l_43 [399] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7079]    = ( l_43 [400] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7080]    = ( l_43 [401] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7081]    = ( l_43 [402] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7082]    = ( l_43 [399] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7083]    = ( l_43 [400] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7084]    = ( l_43 [401] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7085]    = ( l_43 [402] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7086]    = ( l_43 [399] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7087]    = ( l_43 [400] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7088]    = ( l_43 [401] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7089]    = ( l_43 [402] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7090]    = ( l_43 [403] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7091]    = ( l_43 [404] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7092]    = ( l_43 [405] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7093]    = ( l_43 [406] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7094]    = ( l_43 [403] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7095]    = ( l_43 [404] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7096]    = ( l_43 [405] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7097]    = ( l_43 [406] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7098]    = ( l_43 [403] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7099]    = ( l_43 [404] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7100]    = ( l_43 [405] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7101]    = ( l_43 [406] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7102]    = ( l_43 [403] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7103]    = ( l_43 [404] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7104]    = ( l_43 [405] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7105]    = ( l_43 [406] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7106]    = ( l_43 [407] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7107]    = ( l_43 [408] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7108]    = ( l_43 [409] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7109]    = ( l_43 [410] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7110]    = ( l_43 [407] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7111]    = ( l_43 [408] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7112]    = ( l_43 [409] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7113]    = ( l_43 [410] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7114]    = ( l_43 [407] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7115]    = ( l_43 [408] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7116]    = ( l_43 [409] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7117]    = ( l_43 [410] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7118]    = ( l_43 [407] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7119]    = ( l_43 [408] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7120]    = ( l_43 [409] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7121]    = ( l_43 [410] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7122]    = ( l_43 [411] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7123]    = ( l_43 [412] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7124]    = ( l_43 [413] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7125]    = ( l_43 [414] & !i[1703]) | ( l_43 [210] &  i[1703]);
assign l_42[7126]    = ( l_43 [411] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7127]    = ( l_43 [412] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7128]    = ( l_43 [413] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7129]    = ( l_43 [414] & !i[1703]) | ( l_43 [242] &  i[1703]);
assign l_42[7130]    = ( l_43 [411] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7131]    = ( l_43 [412] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7132]    = ( l_43 [413] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7133]    = ( l_43 [414] & !i[1703]) | ( l_43 [211] &  i[1703]);
assign l_42[7134]    = ( l_43 [411] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7135]    = ( l_43 [412] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7136]    = ( l_43 [413] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7137]    = ( l_43 [414] & !i[1703]) | ( l_43 [243] &  i[1703]);
assign l_42[7138]    = ( l_43 [407] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7139]    = ( l_43 [408] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7140]    = ( l_43 [409] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7141]    = ( l_43 [410] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7142]    = ( l_43 [407] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7143]    = ( l_43 [408] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7144]    = ( l_43 [409] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7145]    = ( l_43 [410] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7146]    = ( l_43 [407] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7147]    = ( l_43 [408] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7148]    = ( l_43 [409] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7149]    = ( l_43 [410] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7150]    = ( l_43 [407] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7151]    = ( l_43 [408] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7152]    = ( l_43 [409] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7153]    = ( l_43 [410] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7154]    = ( l_43 [411] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7155]    = ( l_43 [412] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7156]    = ( l_43 [413] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7157]    = ( l_43 [414] & !i[1703]) | ( l_43 [226] &  i[1703]);
assign l_42[7158]    = ( l_43 [411] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7159]    = ( l_43 [412] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7160]    = ( l_43 [413] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7161]    = ( l_43 [414] & !i[1703]) | ( l_43 [258] &  i[1703]);
assign l_42[7162]    = ( l_43 [411] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7163]    = ( l_43 [412] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7164]    = ( l_43 [413] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7165]    = ( l_43 [414] & !i[1703]) | ( l_43 [227] &  i[1703]);
assign l_42[7166]    = ( l_43 [411] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7167]    = ( l_43 [412] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7168]    = ( l_43 [413] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7169]    = ( l_43 [414] & !i[1703]) | ( l_43 [259] &  i[1703]);
assign l_42[7170]    = ( l_43 [407] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7171]    = ( l_43 [408] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7172]    = ( l_43 [409] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7173]    = ( l_43 [410] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7174]    = ( l_43 [407] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7175]    = ( l_43 [408] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7176]    = ( l_43 [409] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7177]    = ( l_43 [410] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7178]    = ( l_43 [407] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7179]    = ( l_43 [408] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7180]    = ( l_43 [409] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7181]    = ( l_43 [410] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7182]    = ( l_43 [407] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7183]    = ( l_43 [408] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7184]    = ( l_43 [409] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7185]    = ( l_43 [410] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7186]    = ( l_43 [411] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7187]    = ( l_43 [412] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7188]    = ( l_43 [413] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7189]    = ( l_43 [414] & !i[1703]) | ( l_43 [214] &  i[1703]);
assign l_42[7190]    = ( l_43 [411] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7191]    = ( l_43 [412] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7192]    = ( l_43 [413] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7193]    = ( l_43 [414] & !i[1703]) | ( l_43 [246] &  i[1703]);
assign l_42[7194]    = ( l_43 [411] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7195]    = ( l_43 [412] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7196]    = ( l_43 [413] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7197]    = ( l_43 [414] & !i[1703]) | ( l_43 [215] &  i[1703]);
assign l_42[7198]    = ( l_43 [411] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7199]    = ( l_43 [412] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7200]    = ( l_43 [413] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7201]    = ( l_43 [414] & !i[1703]) | ( l_43 [247] &  i[1703]);
assign l_42[7202]    = ( l_43 [407] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7203]    = ( l_43 [408] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7204]    = ( l_43 [409] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7205]    = ( l_43 [410] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7206]    = ( l_43 [407] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7207]    = ( l_43 [408] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7208]    = ( l_43 [409] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7209]    = ( l_43 [410] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7210]    = ( l_43 [407] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7211]    = ( l_43 [408] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7212]    = ( l_43 [409] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7213]    = ( l_43 [410] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7214]    = ( l_43 [407] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7215]    = ( l_43 [408] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7216]    = ( l_43 [409] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7217]    = ( l_43 [410] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7218]    = ( l_43 [411] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7219]    = ( l_43 [412] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7220]    = ( l_43 [413] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7221]    = ( l_43 [414] & !i[1703]) | ( l_43 [230] &  i[1703]);
assign l_42[7222]    = ( l_43 [411] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7223]    = ( l_43 [412] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7224]    = ( l_43 [413] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7225]    = ( l_43 [414] & !i[1703]) | ( l_43 [262] &  i[1703]);
assign l_42[7226]    = ( l_43 [411] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7227]    = ( l_43 [412] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7228]    = ( l_43 [413] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7229]    = ( l_43 [414] & !i[1703]) | ( l_43 [231] &  i[1703]);
assign l_42[7230]    = ( l_43 [411] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7231]    = ( l_43 [412] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7232]    = ( l_43 [413] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7233]    = ( l_43 [414] & !i[1703]) | ( l_43 [263] &  i[1703]);
assign l_42[7234]    = ( l_43 [399] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7235]    = ( l_43 [400] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7236]    = ( l_43 [401] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7237]    = ( l_43 [402] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7238]    = ( l_43 [399] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7239]    = ( l_43 [400] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7240]    = ( l_43 [401] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7241]    = ( l_43 [402] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7242]    = ( l_43 [399] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7243]    = ( l_43 [400] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7244]    = ( l_43 [401] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7245]    = ( l_43 [402] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7246]    = ( l_43 [399] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7247]    = ( l_43 [400] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7248]    = ( l_43 [401] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7249]    = ( l_43 [402] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7250]    = ( l_43 [403] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7251]    = ( l_43 [404] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7252]    = ( l_43 [405] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7253]    = ( l_43 [406] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7254]    = ( l_43 [403] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7255]    = ( l_43 [404] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7256]    = ( l_43 [405] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7257]    = ( l_43 [406] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7258]    = ( l_43 [403] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7259]    = ( l_43 [404] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7260]    = ( l_43 [405] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7261]    = ( l_43 [406] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7262]    = ( l_43 [403] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7263]    = ( l_43 [404] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7264]    = ( l_43 [405] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7265]    = ( l_43 [406] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7266]    = ( l_43 [399] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7267]    = ( l_43 [400] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7268]    = ( l_43 [401] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7269]    = ( l_43 [402] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7270]    = ( l_43 [399] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7271]    = ( l_43 [400] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7272]    = ( l_43 [401] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7273]    = ( l_43 [402] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7274]    = ( l_43 [399] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7275]    = ( l_43 [400] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7276]    = ( l_43 [401] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7277]    = ( l_43 [402] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7278]    = ( l_43 [399] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7279]    = ( l_43 [400] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7280]    = ( l_43 [401] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7281]    = ( l_43 [402] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7282]    = ( l_43 [403] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7283]    = ( l_43 [404] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7284]    = ( l_43 [405] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7285]    = ( l_43 [406] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7286]    = ( l_43 [403] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7287]    = ( l_43 [404] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7288]    = ( l_43 [405] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7289]    = ( l_43 [406] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7290]    = ( l_43 [403] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7291]    = ( l_43 [404] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7292]    = ( l_43 [405] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7293]    = ( l_43 [406] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7294]    = ( l_43 [403] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7295]    = ( l_43 [404] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7296]    = ( l_43 [405] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7297]    = ( l_43 [406] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7298]    = ( l_43 [399] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7299]    = ( l_43 [400] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7300]    = ( l_43 [401] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7301]    = ( l_43 [402] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7302]    = ( l_43 [399] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7303]    = ( l_43 [400] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7304]    = ( l_43 [401] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7305]    = ( l_43 [402] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7306]    = ( l_43 [399] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7307]    = ( l_43 [400] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7308]    = ( l_43 [401] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7309]    = ( l_43 [402] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7310]    = ( l_43 [399] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7311]    = ( l_43 [400] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7312]    = ( l_43 [401] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7313]    = ( l_43 [402] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7314]    = ( l_43 [403] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7315]    = ( l_43 [404] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7316]    = ( l_43 [405] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7317]    = ( l_43 [406] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7318]    = ( l_43 [403] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7319]    = ( l_43 [404] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7320]    = ( l_43 [405] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7321]    = ( l_43 [406] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7322]    = ( l_43 [403] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7323]    = ( l_43 [404] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7324]    = ( l_43 [405] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7325]    = ( l_43 [406] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7326]    = ( l_43 [403] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7327]    = ( l_43 [404] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7328]    = ( l_43 [405] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7329]    = ( l_43 [406] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7330]    = ( l_43 [399] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7331]    = ( l_43 [400] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7332]    = ( l_43 [401] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7333]    = ( l_43 [402] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7334]    = ( l_43 [399] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7335]    = ( l_43 [400] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7336]    = ( l_43 [401] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7337]    = ( l_43 [402] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7338]    = ( l_43 [399] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7339]    = ( l_43 [400] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7340]    = ( l_43 [401] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7341]    = ( l_43 [402] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7342]    = ( l_43 [399] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7343]    = ( l_43 [400] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7344]    = ( l_43 [401] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7345]    = ( l_43 [402] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7346]    = ( l_43 [403] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7347]    = ( l_43 [404] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7348]    = ( l_43 [405] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7349]    = ( l_43 [406] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7350]    = ( l_43 [403] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7351]    = ( l_43 [404] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7352]    = ( l_43 [405] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7353]    = ( l_43 [406] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7354]    = ( l_43 [403] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7355]    = ( l_43 [404] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7356]    = ( l_43 [405] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7357]    = ( l_43 [406] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7358]    = ( l_43 [403] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7359]    = ( l_43 [404] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7360]    = ( l_43 [405] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7361]    = ( l_43 [406] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7362]    = ( l_43 [407] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7363]    = ( l_43 [408] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7364]    = ( l_43 [409] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7365]    = ( l_43 [410] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7366]    = ( l_43 [407] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7367]    = ( l_43 [408] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7368]    = ( l_43 [409] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7369]    = ( l_43 [410] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7370]    = ( l_43 [407] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7371]    = ( l_43 [408] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7372]    = ( l_43 [409] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7373]    = ( l_43 [410] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7374]    = ( l_43 [407] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7375]    = ( l_43 [408] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7376]    = ( l_43 [409] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7377]    = ( l_43 [410] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7378]    = ( l_43 [411] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7379]    = ( l_43 [412] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7380]    = ( l_43 [413] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7381]    = ( l_43 [414] & !i[1703]) | ( l_43 [272] &  i[1703]);
assign l_42[7382]    = ( l_43 [411] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7383]    = ( l_43 [412] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7384]    = ( l_43 [413] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7385]    = ( l_43 [414] & !i[1703]) | ( l_43 [304] &  i[1703]);
assign l_42[7386]    = ( l_43 [411] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7387]    = ( l_43 [412] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7388]    = ( l_43 [413] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7389]    = ( l_43 [414] & !i[1703]) | ( l_43 [273] &  i[1703]);
assign l_42[7390]    = ( l_43 [411] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7391]    = ( l_43 [412] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7392]    = ( l_43 [413] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7393]    = ( l_43 [414] & !i[1703]) | ( l_43 [305] &  i[1703]);
assign l_42[7394]    = ( l_43 [407] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7395]    = ( l_43 [408] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7396]    = ( l_43 [409] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7397]    = ( l_43 [410] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7398]    = ( l_43 [407] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7399]    = ( l_43 [408] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7400]    = ( l_43 [409] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7401]    = ( l_43 [410] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7402]    = ( l_43 [407] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7403]    = ( l_43 [408] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7404]    = ( l_43 [409] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7405]    = ( l_43 [410] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7406]    = ( l_43 [407] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7407]    = ( l_43 [408] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7408]    = ( l_43 [409] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7409]    = ( l_43 [410] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7410]    = ( l_43 [411] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7411]    = ( l_43 [412] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7412]    = ( l_43 [413] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7413]    = ( l_43 [414] & !i[1703]) | ( l_43 [288] &  i[1703]);
assign l_42[7414]    = ( l_43 [411] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7415]    = ( l_43 [412] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7416]    = ( l_43 [413] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7417]    = ( l_43 [414] & !i[1703]) | ( l_43 [320] &  i[1703]);
assign l_42[7418]    = ( l_43 [411] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7419]    = ( l_43 [412] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7420]    = ( l_43 [413] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7421]    = ( l_43 [414] & !i[1703]) | ( l_43 [289] &  i[1703]);
assign l_42[7422]    = ( l_43 [411] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7423]    = ( l_43 [412] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7424]    = ( l_43 [413] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7425]    = ( l_43 [414] & !i[1703]) | ( l_43 [321] &  i[1703]);
assign l_42[7426]    = ( l_43 [407] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7427]    = ( l_43 [408] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7428]    = ( l_43 [409] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7429]    = ( l_43 [410] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7430]    = ( l_43 [407] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7431]    = ( l_43 [408] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7432]    = ( l_43 [409] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7433]    = ( l_43 [410] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7434]    = ( l_43 [407] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7435]    = ( l_43 [408] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7436]    = ( l_43 [409] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7437]    = ( l_43 [410] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7438]    = ( l_43 [407] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7439]    = ( l_43 [408] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7440]    = ( l_43 [409] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7441]    = ( l_43 [410] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7442]    = ( l_43 [411] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7443]    = ( l_43 [412] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7444]    = ( l_43 [413] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7445]    = ( l_43 [414] & !i[1703]) | ( l_43 [276] &  i[1703]);
assign l_42[7446]    = ( l_43 [411] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7447]    = ( l_43 [412] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7448]    = ( l_43 [413] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7449]    = ( l_43 [414] & !i[1703]) | ( l_43 [308] &  i[1703]);
assign l_42[7450]    = ( l_43 [411] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7451]    = ( l_43 [412] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7452]    = ( l_43 [413] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7453]    = ( l_43 [414] & !i[1703]) | ( l_43 [277] &  i[1703]);
assign l_42[7454]    = ( l_43 [411] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7455]    = ( l_43 [412] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7456]    = ( l_43 [413] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7457]    = ( l_43 [414] & !i[1703]) | ( l_43 [309] &  i[1703]);
assign l_42[7458]    = ( l_43 [407] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7459]    = ( l_43 [408] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7460]    = ( l_43 [409] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7461]    = ( l_43 [410] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7462]    = ( l_43 [407] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7463]    = ( l_43 [408] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7464]    = ( l_43 [409] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7465]    = ( l_43 [410] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7466]    = ( l_43 [407] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7467]    = ( l_43 [408] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7468]    = ( l_43 [409] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7469]    = ( l_43 [410] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7470]    = ( l_43 [407] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7471]    = ( l_43 [408] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7472]    = ( l_43 [409] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7473]    = ( l_43 [410] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7474]    = ( l_43 [411] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7475]    = ( l_43 [412] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7476]    = ( l_43 [413] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7477]    = ( l_43 [414] & !i[1703]) | ( l_43 [292] &  i[1703]);
assign l_42[7478]    = ( l_43 [411] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7479]    = ( l_43 [412] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7480]    = ( l_43 [413] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7481]    = ( l_43 [414] & !i[1703]) | ( l_43 [324] &  i[1703]);
assign l_42[7482]    = ( l_43 [411] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7483]    = ( l_43 [412] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7484]    = ( l_43 [413] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7485]    = ( l_43 [414] & !i[1703]) | ( l_43 [293] &  i[1703]);
assign l_42[7486]    = ( l_43 [411] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7487]    = ( l_43 [412] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7488]    = ( l_43 [413] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7489]    = ( l_43 [414] & !i[1703]) | ( l_43 [325] &  i[1703]);
assign l_42[7490]    = ( l_43 [399] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7491]    = ( l_43 [400] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7492]    = ( l_43 [401] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7493]    = ( l_43 [402] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7494]    = ( l_43 [399] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7495]    = ( l_43 [400] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7496]    = ( l_43 [401] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7497]    = ( l_43 [402] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7498]    = ( l_43 [399] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7499]    = ( l_43 [400] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7500]    = ( l_43 [401] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7501]    = ( l_43 [402] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7502]    = ( l_43 [399] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7503]    = ( l_43 [400] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7504]    = ( l_43 [401] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7505]    = ( l_43 [402] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7506]    = ( l_43 [403] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7507]    = ( l_43 [404] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7508]    = ( l_43 [405] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7509]    = ( l_43 [406] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7510]    = ( l_43 [403] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7511]    = ( l_43 [404] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7512]    = ( l_43 [405] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7513]    = ( l_43 [406] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7514]    = ( l_43 [403] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7515]    = ( l_43 [404] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7516]    = ( l_43 [405] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7517]    = ( l_43 [406] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7518]    = ( l_43 [403] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7519]    = ( l_43 [404] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7520]    = ( l_43 [405] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7521]    = ( l_43 [406] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7522]    = ( l_43 [399] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7523]    = ( l_43 [400] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7524]    = ( l_43 [401] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7525]    = ( l_43 [402] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7526]    = ( l_43 [399] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7527]    = ( l_43 [400] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7528]    = ( l_43 [401] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7529]    = ( l_43 [402] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7530]    = ( l_43 [399] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7531]    = ( l_43 [400] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7532]    = ( l_43 [401] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7533]    = ( l_43 [402] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7534]    = ( l_43 [399] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7535]    = ( l_43 [400] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7536]    = ( l_43 [401] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7537]    = ( l_43 [402] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7538]    = ( l_43 [403] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7539]    = ( l_43 [404] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7540]    = ( l_43 [405] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7541]    = ( l_43 [406] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7542]    = ( l_43 [403] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7543]    = ( l_43 [404] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7544]    = ( l_43 [405] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7545]    = ( l_43 [406] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7546]    = ( l_43 [403] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7547]    = ( l_43 [404] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7548]    = ( l_43 [405] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7549]    = ( l_43 [406] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7550]    = ( l_43 [403] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7551]    = ( l_43 [404] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7552]    = ( l_43 [405] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7553]    = ( l_43 [406] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7554]    = ( l_43 [399] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7555]    = ( l_43 [400] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7556]    = ( l_43 [401] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7557]    = ( l_43 [402] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7558]    = ( l_43 [399] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7559]    = ( l_43 [400] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7560]    = ( l_43 [401] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7561]    = ( l_43 [402] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7562]    = ( l_43 [399] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7563]    = ( l_43 [400] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7564]    = ( l_43 [401] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7565]    = ( l_43 [402] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7566]    = ( l_43 [399] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7567]    = ( l_43 [400] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7568]    = ( l_43 [401] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7569]    = ( l_43 [402] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7570]    = ( l_43 [403] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7571]    = ( l_43 [404] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7572]    = ( l_43 [405] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7573]    = ( l_43 [406] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7574]    = ( l_43 [403] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7575]    = ( l_43 [404] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7576]    = ( l_43 [405] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7577]    = ( l_43 [406] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7578]    = ( l_43 [403] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7579]    = ( l_43 [404] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7580]    = ( l_43 [405] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7581]    = ( l_43 [406] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7582]    = ( l_43 [403] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7583]    = ( l_43 [404] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7584]    = ( l_43 [405] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7585]    = ( l_43 [406] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7586]    = ( l_43 [399] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7587]    = ( l_43 [400] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7588]    = ( l_43 [401] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7589]    = ( l_43 [402] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7590]    = ( l_43 [399] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7591]    = ( l_43 [400] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7592]    = ( l_43 [401] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7593]    = ( l_43 [402] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7594]    = ( l_43 [399] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7595]    = ( l_43 [400] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7596]    = ( l_43 [401] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7597]    = ( l_43 [402] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7598]    = ( l_43 [399] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7599]    = ( l_43 [400] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7600]    = ( l_43 [401] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7601]    = ( l_43 [402] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7602]    = ( l_43 [403] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7603]    = ( l_43 [404] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7604]    = ( l_43 [405] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7605]    = ( l_43 [406] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7606]    = ( l_43 [403] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7607]    = ( l_43 [404] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7608]    = ( l_43 [405] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7609]    = ( l_43 [406] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7610]    = ( l_43 [403] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7611]    = ( l_43 [404] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7612]    = ( l_43 [405] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7613]    = ( l_43 [406] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7614]    = ( l_43 [403] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7615]    = ( l_43 [404] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7616]    = ( l_43 [405] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7617]    = ( l_43 [406] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7618]    = ( l_43 [407] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7619]    = ( l_43 [408] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7620]    = ( l_43 [409] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7621]    = ( l_43 [410] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7622]    = ( l_43 [407] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7623]    = ( l_43 [408] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7624]    = ( l_43 [409] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7625]    = ( l_43 [410] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7626]    = ( l_43 [407] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7627]    = ( l_43 [408] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7628]    = ( l_43 [409] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7629]    = ( l_43 [410] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7630]    = ( l_43 [407] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7631]    = ( l_43 [408] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7632]    = ( l_43 [409] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7633]    = ( l_43 [410] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7634]    = ( l_43 [411] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7635]    = ( l_43 [412] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7636]    = ( l_43 [413] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7637]    = ( l_43 [414] & !i[1703]) | ( l_43 [274] &  i[1703]);
assign l_42[7638]    = ( l_43 [411] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7639]    = ( l_43 [412] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7640]    = ( l_43 [413] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7641]    = ( l_43 [414] & !i[1703]) | ( l_43 [306] &  i[1703]);
assign l_42[7642]    = ( l_43 [411] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7643]    = ( l_43 [412] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7644]    = ( l_43 [413] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7645]    = ( l_43 [414] & !i[1703]) | ( l_43 [275] &  i[1703]);
assign l_42[7646]    = ( l_43 [411] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7647]    = ( l_43 [412] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7648]    = ( l_43 [413] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7649]    = ( l_43 [414] & !i[1703]) | ( l_43 [307] &  i[1703]);
assign l_42[7650]    = ( l_43 [407] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7651]    = ( l_43 [408] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7652]    = ( l_43 [409] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7653]    = ( l_43 [410] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7654]    = ( l_43 [407] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7655]    = ( l_43 [408] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7656]    = ( l_43 [409] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7657]    = ( l_43 [410] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7658]    = ( l_43 [407] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7659]    = ( l_43 [408] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7660]    = ( l_43 [409] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7661]    = ( l_43 [410] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7662]    = ( l_43 [407] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7663]    = ( l_43 [408] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7664]    = ( l_43 [409] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7665]    = ( l_43 [410] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7666]    = ( l_43 [411] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7667]    = ( l_43 [412] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7668]    = ( l_43 [413] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7669]    = ( l_43 [414] & !i[1703]) | ( l_43 [290] &  i[1703]);
assign l_42[7670]    = ( l_43 [411] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7671]    = ( l_43 [412] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7672]    = ( l_43 [413] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7673]    = ( l_43 [414] & !i[1703]) | ( l_43 [322] &  i[1703]);
assign l_42[7674]    = ( l_43 [411] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7675]    = ( l_43 [412] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7676]    = ( l_43 [413] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7677]    = ( l_43 [414] & !i[1703]) | ( l_43 [291] &  i[1703]);
assign l_42[7678]    = ( l_43 [411] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7679]    = ( l_43 [412] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7680]    = ( l_43 [413] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7681]    = ( l_43 [414] & !i[1703]) | ( l_43 [323] &  i[1703]);
assign l_42[7682]    = ( l_43 [407] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7683]    = ( l_43 [408] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7684]    = ( l_43 [409] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7685]    = ( l_43 [410] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7686]    = ( l_43 [407] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7687]    = ( l_43 [408] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7688]    = ( l_43 [409] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7689]    = ( l_43 [410] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7690]    = ( l_43 [407] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7691]    = ( l_43 [408] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7692]    = ( l_43 [409] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7693]    = ( l_43 [410] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7694]    = ( l_43 [407] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7695]    = ( l_43 [408] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7696]    = ( l_43 [409] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7697]    = ( l_43 [410] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7698]    = ( l_43 [411] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7699]    = ( l_43 [412] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7700]    = ( l_43 [413] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7701]    = ( l_43 [414] & !i[1703]) | ( l_43 [278] &  i[1703]);
assign l_42[7702]    = ( l_43 [411] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7703]    = ( l_43 [412] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7704]    = ( l_43 [413] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7705]    = ( l_43 [414] & !i[1703]) | ( l_43 [310] &  i[1703]);
assign l_42[7706]    = ( l_43 [411] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7707]    = ( l_43 [412] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7708]    = ( l_43 [413] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7709]    = ( l_43 [414] & !i[1703]) | ( l_43 [279] &  i[1703]);
assign l_42[7710]    = ( l_43 [411] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7711]    = ( l_43 [412] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7712]    = ( l_43 [413] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7713]    = ( l_43 [414] & !i[1703]) | ( l_43 [311] &  i[1703]);
assign l_42[7714]    = ( l_43 [407] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7715]    = ( l_43 [408] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7716]    = ( l_43 [409] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7717]    = ( l_43 [410] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7718]    = ( l_43 [407] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7719]    = ( l_43 [408] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7720]    = ( l_43 [409] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7721]    = ( l_43 [410] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7722]    = ( l_43 [407] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7723]    = ( l_43 [408] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7724]    = ( l_43 [409] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7725]    = ( l_43 [410] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7726]    = ( l_43 [407] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7727]    = ( l_43 [408] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7728]    = ( l_43 [409] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7729]    = ( l_43 [410] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7730]    = ( l_43 [411] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7731]    = ( l_43 [412] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7732]    = ( l_43 [413] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7733]    = ( l_43 [414] & !i[1703]) | ( l_43 [294] &  i[1703]);
assign l_42[7734]    = ( l_43 [411] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7735]    = ( l_43 [412] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7736]    = ( l_43 [413] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7737]    = ( l_43 [414] & !i[1703]) | ( l_43 [326] &  i[1703]);
assign l_42[7738]    = ( l_43 [411] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7739]    = ( l_43 [412] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7740]    = ( l_43 [413] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7741]    = ( l_43 [414] & !i[1703]) | ( l_43 [295] &  i[1703]);
assign l_42[7742]    = ( l_43 [411] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7743]    = ( l_43 [412] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7744]    = ( l_43 [413] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7745]    = ( l_43 [414] & !i[1703]) | ( l_43 [327] &  i[1703]);
assign l_42[7746]    = ( l_43 [399] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7747]    = ( l_43 [400] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7748]    = ( l_43 [401] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7749]    = ( l_43 [402] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7750]    = ( l_43 [399] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7751]    = ( l_43 [400] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7752]    = ( l_43 [401] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7753]    = ( l_43 [402] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7754]    = ( l_43 [399] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7755]    = ( l_43 [400] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7756]    = ( l_43 [401] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7757]    = ( l_43 [402] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7758]    = ( l_43 [399] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7759]    = ( l_43 [400] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7760]    = ( l_43 [401] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7761]    = ( l_43 [402] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7762]    = ( l_43 [403] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7763]    = ( l_43 [404] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7764]    = ( l_43 [405] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7765]    = ( l_43 [406] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7766]    = ( l_43 [403] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7767]    = ( l_43 [404] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7768]    = ( l_43 [405] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7769]    = ( l_43 [406] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7770]    = ( l_43 [403] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7771]    = ( l_43 [404] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7772]    = ( l_43 [405] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7773]    = ( l_43 [406] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7774]    = ( l_43 [403] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7775]    = ( l_43 [404] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7776]    = ( l_43 [405] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7777]    = ( l_43 [406] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7778]    = ( l_43 [399] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7779]    = ( l_43 [400] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7780]    = ( l_43 [401] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7781]    = ( l_43 [402] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7782]    = ( l_43 [399] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7783]    = ( l_43 [400] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7784]    = ( l_43 [401] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7785]    = ( l_43 [402] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7786]    = ( l_43 [399] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7787]    = ( l_43 [400] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7788]    = ( l_43 [401] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7789]    = ( l_43 [402] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7790]    = ( l_43 [399] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7791]    = ( l_43 [400] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7792]    = ( l_43 [401] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7793]    = ( l_43 [402] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7794]    = ( l_43 [403] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7795]    = ( l_43 [404] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7796]    = ( l_43 [405] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7797]    = ( l_43 [406] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7798]    = ( l_43 [403] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7799]    = ( l_43 [404] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7800]    = ( l_43 [405] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7801]    = ( l_43 [406] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7802]    = ( l_43 [403] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7803]    = ( l_43 [404] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7804]    = ( l_43 [405] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7805]    = ( l_43 [406] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7806]    = ( l_43 [403] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7807]    = ( l_43 [404] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7808]    = ( l_43 [405] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7809]    = ( l_43 [406] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7810]    = ( l_43 [399] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7811]    = ( l_43 [400] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7812]    = ( l_43 [401] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7813]    = ( l_43 [402] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7814]    = ( l_43 [399] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7815]    = ( l_43 [400] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7816]    = ( l_43 [401] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7817]    = ( l_43 [402] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7818]    = ( l_43 [399] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7819]    = ( l_43 [400] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7820]    = ( l_43 [401] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7821]    = ( l_43 [402] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7822]    = ( l_43 [399] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7823]    = ( l_43 [400] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7824]    = ( l_43 [401] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7825]    = ( l_43 [402] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7826]    = ( l_43 [403] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7827]    = ( l_43 [404] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7828]    = ( l_43 [405] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7829]    = ( l_43 [406] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7830]    = ( l_43 [403] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7831]    = ( l_43 [404] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7832]    = ( l_43 [405] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7833]    = ( l_43 [406] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7834]    = ( l_43 [403] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7835]    = ( l_43 [404] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7836]    = ( l_43 [405] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7837]    = ( l_43 [406] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7838]    = ( l_43 [403] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7839]    = ( l_43 [404] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7840]    = ( l_43 [405] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7841]    = ( l_43 [406] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7842]    = ( l_43 [399] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7843]    = ( l_43 [400] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7844]    = ( l_43 [401] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7845]    = ( l_43 [402] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7846]    = ( l_43 [399] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7847]    = ( l_43 [400] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7848]    = ( l_43 [401] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7849]    = ( l_43 [402] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7850]    = ( l_43 [399] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7851]    = ( l_43 [400] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7852]    = ( l_43 [401] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7853]    = ( l_43 [402] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7854]    = ( l_43 [399] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7855]    = ( l_43 [400] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7856]    = ( l_43 [401] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7857]    = ( l_43 [402] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7858]    = ( l_43 [403] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7859]    = ( l_43 [404] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7860]    = ( l_43 [405] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7861]    = ( l_43 [406] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7862]    = ( l_43 [403] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7863]    = ( l_43 [404] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7864]    = ( l_43 [405] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7865]    = ( l_43 [406] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7866]    = ( l_43 [403] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7867]    = ( l_43 [404] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7868]    = ( l_43 [405] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7869]    = ( l_43 [406] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7870]    = ( l_43 [403] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7871]    = ( l_43 [404] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7872]    = ( l_43 [405] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7873]    = ( l_43 [406] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7874]    = ( l_43 [407] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7875]    = ( l_43 [408] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7876]    = ( l_43 [409] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7877]    = ( l_43 [410] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7878]    = ( l_43 [407] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7879]    = ( l_43 [408] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7880]    = ( l_43 [409] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7881]    = ( l_43 [410] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7882]    = ( l_43 [407] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7883]    = ( l_43 [408] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7884]    = ( l_43 [409] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7885]    = ( l_43 [410] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7886]    = ( l_43 [407] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7887]    = ( l_43 [408] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7888]    = ( l_43 [409] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7889]    = ( l_43 [410] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7890]    = ( l_43 [411] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7891]    = ( l_43 [412] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7892]    = ( l_43 [413] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7893]    = ( l_43 [414] & !i[1703]) | ( l_43 [336] &  i[1703]);
assign l_42[7894]    = ( l_43 [411] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7895]    = ( l_43 [412] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7896]    = ( l_43 [413] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7897]    = ( l_43 [414] & !i[1703]) | ( l_43 [368] &  i[1703]);
assign l_42[7898]    = ( l_43 [411] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7899]    = ( l_43 [412] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7900]    = ( l_43 [413] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7901]    = ( l_43 [414] & !i[1703]) | ( l_43 [337] &  i[1703]);
assign l_42[7902]    = ( l_43 [411] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7903]    = ( l_43 [412] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7904]    = ( l_43 [413] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7905]    = ( l_43 [414] & !i[1703]) | ( l_43 [369] &  i[1703]);
assign l_42[7906]    = ( l_43 [407] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7907]    = ( l_43 [408] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7908]    = ( l_43 [409] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7909]    = ( l_43 [410] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7910]    = ( l_43 [407] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7911]    = ( l_43 [408] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7912]    = ( l_43 [409] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7913]    = ( l_43 [410] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7914]    = ( l_43 [407] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7915]    = ( l_43 [408] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7916]    = ( l_43 [409] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7917]    = ( l_43 [410] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7918]    = ( l_43 [407] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7919]    = ( l_43 [408] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7920]    = ( l_43 [409] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7921]    = ( l_43 [410] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7922]    = ( l_43 [411] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7923]    = ( l_43 [412] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7924]    = ( l_43 [413] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7925]    = ( l_43 [414] & !i[1703]) | ( l_43 [352] &  i[1703]);
assign l_42[7926]    = ( l_43 [411] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7927]    = ( l_43 [412] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7928]    = ( l_43 [413] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7929]    = ( l_43 [414] & !i[1703]) | ( l_43 [384] &  i[1703]);
assign l_42[7930]    = ( l_43 [411] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7931]    = ( l_43 [412] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7932]    = ( l_43 [413] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7933]    = ( l_43 [414] & !i[1703]) | ( l_43 [353] &  i[1703]);
assign l_42[7934]    = ( l_43 [411] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7935]    = ( l_43 [412] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7936]    = ( l_43 [413] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7937]    = ( l_43 [414] & !i[1703]) | ( l_43 [385] &  i[1703]);
assign l_42[7938]    = ( l_43 [407] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7939]    = ( l_43 [408] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7940]    = ( l_43 [409] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7941]    = ( l_43 [410] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7942]    = ( l_43 [407] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7943]    = ( l_43 [408] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7944]    = ( l_43 [409] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7945]    = ( l_43 [410] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7946]    = ( l_43 [407] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7947]    = ( l_43 [408] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7948]    = ( l_43 [409] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7949]    = ( l_43 [410] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7950]    = ( l_43 [407] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7951]    = ( l_43 [408] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7952]    = ( l_43 [409] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7953]    = ( l_43 [410] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7954]    = ( l_43 [411] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7955]    = ( l_43 [412] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7956]    = ( l_43 [413] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7957]    = ( l_43 [414] & !i[1703]) | ( l_43 [340] &  i[1703]);
assign l_42[7958]    = ( l_43 [411] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7959]    = ( l_43 [412] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7960]    = ( l_43 [413] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7961]    = ( l_43 [414] & !i[1703]) | ( l_43 [372] &  i[1703]);
assign l_42[7962]    = ( l_43 [411] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7963]    = ( l_43 [412] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7964]    = ( l_43 [413] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7965]    = ( l_43 [414] & !i[1703]) | ( l_43 [341] &  i[1703]);
assign l_42[7966]    = ( l_43 [411] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7967]    = ( l_43 [412] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7968]    = ( l_43 [413] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7969]    = ( l_43 [414] & !i[1703]) | ( l_43 [373] &  i[1703]);
assign l_42[7970]    = ( l_43 [407] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7971]    = ( l_43 [408] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7972]    = ( l_43 [409] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7973]    = ( l_43 [410] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7974]    = ( l_43 [407] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7975]    = ( l_43 [408] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7976]    = ( l_43 [409] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7977]    = ( l_43 [410] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7978]    = ( l_43 [407] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7979]    = ( l_43 [408] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7980]    = ( l_43 [409] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7981]    = ( l_43 [410] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7982]    = ( l_43 [407] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7983]    = ( l_43 [408] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7984]    = ( l_43 [409] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7985]    = ( l_43 [410] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7986]    = ( l_43 [411] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7987]    = ( l_43 [412] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7988]    = ( l_43 [413] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7989]    = ( l_43 [414] & !i[1703]) | ( l_43 [356] &  i[1703]);
assign l_42[7990]    = ( l_43 [411] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7991]    = ( l_43 [412] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7992]    = ( l_43 [413] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7993]    = ( l_43 [414] & !i[1703]) | ( l_43 [388] &  i[1703]);
assign l_42[7994]    = ( l_43 [411] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7995]    = ( l_43 [412] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7996]    = ( l_43 [413] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7997]    = ( l_43 [414] & !i[1703]) | ( l_43 [357] &  i[1703]);
assign l_42[7998]    = ( l_43 [411] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[7999]    = ( l_43 [412] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[8000]    = ( l_43 [413] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[8001]    = ( l_43 [414] & !i[1703]) | ( l_43 [389] &  i[1703]);
assign l_42[8002]    = ( l_43 [399] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8003]    = ( l_43 [400] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8004]    = ( l_43 [401] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8005]    = ( l_43 [402] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8006]    = ( l_43 [399] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8007]    = ( l_43 [400] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8008]    = ( l_43 [401] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8009]    = ( l_43 [402] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8010]    = ( l_43 [399] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8011]    = ( l_43 [400] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8012]    = ( l_43 [401] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8013]    = ( l_43 [402] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8014]    = ( l_43 [399] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8015]    = ( l_43 [400] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8016]    = ( l_43 [401] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8017]    = ( l_43 [402] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8018]    = ( l_43 [403] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8019]    = ( l_43 [404] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8020]    = ( l_43 [405] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8021]    = ( l_43 [406] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8022]    = ( l_43 [403] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8023]    = ( l_43 [404] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8024]    = ( l_43 [405] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8025]    = ( l_43 [406] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8026]    = ( l_43 [403] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8027]    = ( l_43 [404] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8028]    = ( l_43 [405] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8029]    = ( l_43 [406] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8030]    = ( l_43 [403] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8031]    = ( l_43 [404] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8032]    = ( l_43 [405] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8033]    = ( l_43 [406] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8034]    = ( l_43 [399] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8035]    = ( l_43 [400] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8036]    = ( l_43 [401] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8037]    = ( l_43 [402] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8038]    = ( l_43 [399] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8039]    = ( l_43 [400] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8040]    = ( l_43 [401] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8041]    = ( l_43 [402] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8042]    = ( l_43 [399] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8043]    = ( l_43 [400] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8044]    = ( l_43 [401] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8045]    = ( l_43 [402] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8046]    = ( l_43 [399] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8047]    = ( l_43 [400] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8048]    = ( l_43 [401] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8049]    = ( l_43 [402] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8050]    = ( l_43 [403] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8051]    = ( l_43 [404] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8052]    = ( l_43 [405] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8053]    = ( l_43 [406] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8054]    = ( l_43 [403] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8055]    = ( l_43 [404] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8056]    = ( l_43 [405] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8057]    = ( l_43 [406] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8058]    = ( l_43 [403] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8059]    = ( l_43 [404] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8060]    = ( l_43 [405] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8061]    = ( l_43 [406] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8062]    = ( l_43 [403] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8063]    = ( l_43 [404] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8064]    = ( l_43 [405] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8065]    = ( l_43 [406] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8066]    = ( l_43 [399] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8067]    = ( l_43 [400] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8068]    = ( l_43 [401] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8069]    = ( l_43 [402] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8070]    = ( l_43 [399] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8071]    = ( l_43 [400] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8072]    = ( l_43 [401] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8073]    = ( l_43 [402] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8074]    = ( l_43 [399] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8075]    = ( l_43 [400] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8076]    = ( l_43 [401] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8077]    = ( l_43 [402] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8078]    = ( l_43 [399] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8079]    = ( l_43 [400] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8080]    = ( l_43 [401] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8081]    = ( l_43 [402] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8082]    = ( l_43 [403] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8083]    = ( l_43 [404] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8084]    = ( l_43 [405] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8085]    = ( l_43 [406] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8086]    = ( l_43 [403] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8087]    = ( l_43 [404] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8088]    = ( l_43 [405] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8089]    = ( l_43 [406] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8090]    = ( l_43 [403] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8091]    = ( l_43 [404] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8092]    = ( l_43 [405] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8093]    = ( l_43 [406] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8094]    = ( l_43 [403] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8095]    = ( l_43 [404] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8096]    = ( l_43 [405] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8097]    = ( l_43 [406] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8098]    = ( l_43 [399] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8099]    = ( l_43 [400] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8100]    = ( l_43 [401] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8101]    = ( l_43 [402] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8102]    = ( l_43 [399] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8103]    = ( l_43 [400] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8104]    = ( l_43 [401] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8105]    = ( l_43 [402] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8106]    = ( l_43 [399] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8107]    = ( l_43 [400] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8108]    = ( l_43 [401] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8109]    = ( l_43 [402] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8110]    = ( l_43 [399] & !i[1703]) | (      i[1703]);
assign l_42[8111]    = ( l_43 [400] & !i[1703]) | (      i[1703]);
assign l_42[8112]    = ( l_43 [401] & !i[1703]) | (      i[1703]);
assign l_42[8113]    = ( l_43 [402] & !i[1703]) | (      i[1703]);
assign l_42[8114]    = ( l_43 [403] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8115]    = ( l_43 [404] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8116]    = ( l_43 [405] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8117]    = ( l_43 [406] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8118]    = ( l_43 [403] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8119]    = ( l_43 [404] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8120]    = ( l_43 [405] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8121]    = ( l_43 [406] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8122]    = ( l_43 [403] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8123]    = ( l_43 [404] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8124]    = ( l_43 [405] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8125]    = ( l_43 [406] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8126]    = ( l_43 [403] & !i[1703]) | (      i[1703]);
assign l_42[8127]    = ( l_43 [404] & !i[1703]) | (      i[1703]);
assign l_42[8128]    = ( l_43 [405] & !i[1703]) | (      i[1703]);
assign l_42[8129]    = ( l_43 [406] & !i[1703]) | (      i[1703]);
assign l_42[8130]    = ( l_43 [407] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8131]    = ( l_43 [408] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8132]    = ( l_43 [409] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8133]    = ( l_43 [410] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8134]    = ( l_43 [407] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8135]    = ( l_43 [408] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8136]    = ( l_43 [409] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8137]    = ( l_43 [410] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8138]    = ( l_43 [407] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8139]    = ( l_43 [408] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8140]    = ( l_43 [409] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8141]    = ( l_43 [410] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8142]    = ( l_43 [407] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8143]    = ( l_43 [408] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8144]    = ( l_43 [409] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8145]    = ( l_43 [410] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8146]    = ( l_43 [411] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8147]    = ( l_43 [412] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8148]    = ( l_43 [413] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8149]    = ( l_43 [414] & !i[1703]) | ( l_43 [338] &  i[1703]);
assign l_42[8150]    = ( l_43 [411] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8151]    = ( l_43 [412] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8152]    = ( l_43 [413] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8153]    = ( l_43 [414] & !i[1703]) | ( l_43 [370] &  i[1703]);
assign l_42[8154]    = ( l_43 [411] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8155]    = ( l_43 [412] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8156]    = ( l_43 [413] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8157]    = ( l_43 [414] & !i[1703]) | ( l_43 [339] &  i[1703]);
assign l_42[8158]    = ( l_43 [411] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8159]    = ( l_43 [412] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8160]    = ( l_43 [413] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8161]    = ( l_43 [414] & !i[1703]) | ( l_43 [371] &  i[1703]);
assign l_42[8162]    = ( l_43 [407] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8163]    = ( l_43 [408] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8164]    = ( l_43 [409] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8165]    = ( l_43 [410] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8166]    = ( l_43 [407] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8167]    = ( l_43 [408] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8168]    = ( l_43 [409] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8169]    = ( l_43 [410] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8170]    = ( l_43 [407] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8171]    = ( l_43 [408] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8172]    = ( l_43 [409] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8173]    = ( l_43 [410] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8174]    = ( l_43 [407] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8175]    = ( l_43 [408] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8176]    = ( l_43 [409] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8177]    = ( l_43 [410] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8178]    = ( l_43 [411] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8179]    = ( l_43 [412] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8180]    = ( l_43 [413] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8181]    = ( l_43 [414] & !i[1703]) | ( l_43 [354] &  i[1703]);
assign l_42[8182]    = ( l_43 [411] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8183]    = ( l_43 [412] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8184]    = ( l_43 [413] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8185]    = ( l_43 [414] & !i[1703]) | ( l_43 [386] &  i[1703]);
assign l_42[8186]    = ( l_43 [411] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8187]    = ( l_43 [412] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8188]    = ( l_43 [413] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8189]    = ( l_43 [414] & !i[1703]) | ( l_43 [355] &  i[1703]);
assign l_42[8190]    = ( l_43 [411] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8191]    = ( l_43 [412] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8192]    = ( l_43 [413] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8193]    = ( l_43 [414] & !i[1703]) | ( l_43 [387] &  i[1703]);
assign l_42[8194]    = ( l_43 [407] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8195]    = ( l_43 [408] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8196]    = ( l_43 [409] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8197]    = ( l_43 [410] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8198]    = ( l_43 [407] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8199]    = ( l_43 [408] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8200]    = ( l_43 [409] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8201]    = ( l_43 [410] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8202]    = ( l_43 [407] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8203]    = ( l_43 [408] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8204]    = ( l_43 [409] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8205]    = ( l_43 [410] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8206]    = ( l_43 [407] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8207]    = ( l_43 [408] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8208]    = ( l_43 [409] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8209]    = ( l_43 [410] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8210]    = ( l_43 [411] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8211]    = ( l_43 [412] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8212]    = ( l_43 [413] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8213]    = ( l_43 [414] & !i[1703]) | ( l_43 [342] &  i[1703]);
assign l_42[8214]    = ( l_43 [411] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8215]    = ( l_43 [412] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8216]    = ( l_43 [413] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8217]    = ( l_43 [414] & !i[1703]) | ( l_43 [374] &  i[1703]);
assign l_42[8218]    = ( l_43 [411] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8219]    = ( l_43 [412] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8220]    = ( l_43 [413] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8221]    = ( l_43 [414] & !i[1703]) | ( l_43 [343] &  i[1703]);
assign l_42[8222]    = ( l_43 [411] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8223]    = ( l_43 [412] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8224]    = ( l_43 [413] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8225]    = ( l_43 [414] & !i[1703]) | ( l_43 [375] &  i[1703]);
assign l_42[8226]    = ( l_43 [407] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8227]    = ( l_43 [408] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8228]    = ( l_43 [409] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8229]    = ( l_43 [410] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8230]    = ( l_43 [407] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8231]    = ( l_43 [408] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8232]    = ( l_43 [409] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8233]    = ( l_43 [410] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8234]    = ( l_43 [407] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8235]    = ( l_43 [408] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8236]    = ( l_43 [409] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8237]    = ( l_43 [410] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8238]    = ( l_43 [407] & !i[1703]) | (      i[1703]);
assign l_42[8239]    = ( l_43 [408] & !i[1703]) | (      i[1703]);
assign l_42[8240]    = ( l_43 [409] & !i[1703]) | (      i[1703]);
assign l_42[8241]    = ( l_43 [410] & !i[1703]) | (      i[1703]);
assign l_42[8242]    = ( l_43 [411] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8243]    = ( l_43 [412] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8244]    = ( l_43 [413] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8245]    = ( l_43 [414] & !i[1703]) | ( l_43 [358] &  i[1703]);
assign l_42[8246]    = ( l_43 [411] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8247]    = ( l_43 [412] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8248]    = ( l_43 [413] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8249]    = ( l_43 [414] & !i[1703]) | ( l_43 [390] &  i[1703]);
assign l_42[8250]    = ( l_43 [411] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8251]    = ( l_43 [412] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8252]    = ( l_43 [413] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8253]    = ( l_43 [414] & !i[1703]) | ( l_43 [359] &  i[1703]);
assign l_42[8254]    = ( l_43 [411] & !i[1703]) | (      i[1703]);
assign l_42[8255]    = ( l_43 [412] & !i[1703]) | (      i[1703]);
assign l_42[8256]    = ( l_43 [413] & !i[1703]) | (      i[1703]);
assign l_42[8257]    = ( l_43 [414] & !i[1703]) | (      i[1703]);
assign l_43[0]    = ( l_44 [0] & !i[1704]);
assign l_43[1]    = ( l_44 [1] & !i[1704]) | ( l_44 [2] &  i[1704]);
assign l_43[2]    = ( l_44 [3] & !i[1704]) | ( l_44 [4] &  i[1704]);
assign l_43[3]    = ( l_44 [5] & !i[1704]) | ( l_44 [6] &  i[1704]);
assign l_43[4]    = ( l_44 [7] & !i[1704]) | ( l_44 [8] &  i[1704]);
assign l_43[5]    = ( l_44 [9] & !i[1704]) | ( l_44 [10] &  i[1704]);
assign l_43[6]    = ( l_44 [11] & !i[1704]) | ( l_44 [12] &  i[1704]);
assign l_43[7]    = ( l_44 [13] & !i[1704]) | ( l_44 [14] &  i[1704]);
assign l_43[8]    = ( l_44 [15] & !i[1704]) | ( l_44 [16] &  i[1704]);
assign l_43[9]    = ( l_44 [17] & !i[1704]) | ( l_44 [18] &  i[1704]);
assign l_43[10]    = ( l_44 [19] & !i[1704]) | ( l_44 [20] &  i[1704]);
assign l_43[11]    = ( l_44 [21] & !i[1704]) | ( l_44 [22] &  i[1704]);
assign l_43[12]    = ( l_44 [23] & !i[1704]) | ( l_44 [24] &  i[1704]);
assign l_43[13]    = ( l_44 [25] & !i[1704]) | ( l_44 [26] &  i[1704]);
assign l_43[14]    = ( l_44 [27] & !i[1704]) | ( l_44 [28] &  i[1704]);
assign l_43[15]    = ( l_44 [29] & !i[1704]) | ( l_44 [30] &  i[1704]);
assign l_43[16]    = ( l_44 [31] & !i[1704]) | ( l_44 [32] &  i[1704]);
assign l_43[17]    = ( l_44 [33] & !i[1704]) | ( l_44 [34] &  i[1704]);
assign l_43[18]    = ( l_44 [35] & !i[1704]) | ( l_44 [36] &  i[1704]);
assign l_43[19]    = ( l_44 [37] & !i[1704]) | ( l_44 [38] &  i[1704]);
assign l_43[20]    = ( l_44 [39] & !i[1704]) | ( l_44 [40] &  i[1704]);
assign l_43[21]    = ( l_44 [41] & !i[1704]) | ( l_44 [42] &  i[1704]);
assign l_43[22]    = ( l_44 [43] & !i[1704]) | ( l_44 [44] &  i[1704]);
assign l_43[23]    = ( l_44 [45] & !i[1704]) | ( l_44 [46] &  i[1704]);
assign l_43[24]    = ( l_44 [47] & !i[1704]) | ( l_44 [48] &  i[1704]);
assign l_43[25]    = ( l_44 [49] & !i[1704]) | ( l_44 [50] &  i[1704]);
assign l_43[26]    = ( l_44 [51] & !i[1704]) | ( l_44 [52] &  i[1704]);
assign l_43[27]    = ( l_44 [53] & !i[1704]) | ( l_44 [54] &  i[1704]);
assign l_43[28]    = ( l_44 [55] & !i[1704]) | ( l_44 [56] &  i[1704]);
assign l_43[29]    = ( l_44 [57] & !i[1704]) | ( l_44 [58] &  i[1704]);
assign l_43[30]    = ( l_44 [59] & !i[1704]) | ( l_44 [60] &  i[1704]);
assign l_43[31]    = ( l_44 [61] & !i[1704]) | ( l_44 [62] &  i[1704]);
assign l_43[32]    = ( l_44 [63] & !i[1704]) | ( l_44 [64] &  i[1704]);
assign l_43[33]    = ( l_44 [65] & !i[1704]) | ( l_44 [66] &  i[1704]);
assign l_43[34]    = ( l_44 [67] & !i[1704]) | ( l_44 [68] &  i[1704]);
assign l_43[35]    = ( l_44 [69] & !i[1704]) | ( l_44 [70] &  i[1704]);
assign l_43[36]    = ( l_44 [71] & !i[1704]) | ( l_44 [72] &  i[1704]);
assign l_43[37]    = ( l_44 [73] & !i[1704]) | ( l_44 [74] &  i[1704]);
assign l_43[38]    = ( l_44 [75] & !i[1704]) | ( l_44 [76] &  i[1704]);
assign l_43[39]    = ( l_44 [77] & !i[1704]) | ( l_44 [78] &  i[1704]);
assign l_43[40]    = ( l_44 [79] & !i[1704]) | ( l_44 [80] &  i[1704]);
assign l_43[41]    = ( l_44 [81] & !i[1704]) | ( l_44 [82] &  i[1704]);
assign l_43[42]    = ( l_44 [83] & !i[1704]) | ( l_44 [84] &  i[1704]);
assign l_43[43]    = ( l_44 [85] & !i[1704]) | ( l_44 [86] &  i[1704]);
assign l_43[44]    = ( l_44 [87] & !i[1704]) | ( l_44 [88] &  i[1704]);
assign l_43[45]    = ( l_44 [89] & !i[1704]) | ( l_44 [90] &  i[1704]);
assign l_43[46]    = ( l_44 [91] & !i[1704]) | ( l_44 [92] &  i[1704]);
assign l_43[47]    = ( l_44 [93] & !i[1704]) | ( l_44 [94] &  i[1704]);
assign l_43[48]    = ( l_44 [95] & !i[1704]) | ( l_44 [96] &  i[1704]);
assign l_43[49]    = ( l_44 [97] & !i[1704]) | ( l_44 [98] &  i[1704]);
assign l_43[50]    = ( l_44 [99] & !i[1704]) | ( l_44 [100] &  i[1704]);
assign l_43[51]    = ( l_44 [101] & !i[1704]) | ( l_44 [102] &  i[1704]);
assign l_43[52]    = ( l_44 [103] & !i[1704]) | ( l_44 [104] &  i[1704]);
assign l_43[53]    = ( l_44 [105] & !i[1704]) | ( l_44 [106] &  i[1704]);
assign l_43[54]    = ( l_44 [107] & !i[1704]) | ( l_44 [108] &  i[1704]);
assign l_43[55]    = ( l_44 [109] & !i[1704]) | ( l_44 [110] &  i[1704]);
assign l_43[56]    = ( l_44 [111] & !i[1704]) | ( l_44 [112] &  i[1704]);
assign l_43[57]    = ( l_44 [113] & !i[1704]) | ( l_44 [114] &  i[1704]);
assign l_43[58]    = ( l_44 [115] & !i[1704]) | ( l_44 [116] &  i[1704]);
assign l_43[59]    = ( l_44 [117] & !i[1704]) | ( l_44 [118] &  i[1704]);
assign l_43[60]    = ( l_44 [119] & !i[1704]) | ( l_44 [120] &  i[1704]);
assign l_43[61]    = ( l_44 [121] & !i[1704]) | ( l_44 [122] &  i[1704]);
assign l_43[62]    = ( l_44 [123] & !i[1704]) | ( l_44 [124] &  i[1704]);
assign l_43[63]    = ( l_44 [125] & !i[1704]) | ( l_44 [126] &  i[1704]);
assign l_43[64]    = ( l_44 [127] & !i[1704]) | ( l_44 [128] &  i[1704]);
assign l_43[65]    = ( l_44 [129] & !i[1704]) | ( l_44 [130] &  i[1704]);
assign l_43[66]    = ( l_44 [131] & !i[1704]) | ( l_44 [132] &  i[1704]);
assign l_43[67]    = ( l_44 [133] & !i[1704]) | ( l_44 [134] &  i[1704]);
assign l_43[68]    = ( l_44 [135] & !i[1704]) | ( l_44 [136] &  i[1704]);
assign l_43[69]    = ( l_44 [137] & !i[1704]) | ( l_44 [138] &  i[1704]);
assign l_43[70]    = ( l_44 [139] & !i[1704]) | ( l_44 [140] &  i[1704]);
assign l_43[71]    = ( l_44 [141] & !i[1704]) | ( l_44 [142] &  i[1704]);
assign l_43[72]    = ( l_44 [143] & !i[1704]) | ( l_44 [144] &  i[1704]);
assign l_43[73]    = ( l_44 [145]);
assign l_43[74]    = ( l_44 [146] & !i[1704]) | ( l_44 [147] &  i[1704]);
assign l_43[75]    = ( l_44 [148] & !i[1704]) | ( l_44 [149] &  i[1704]);
assign l_43[76]    = ( l_44 [150] & !i[1704]) | ( l_44 [151] &  i[1704]);
assign l_43[77]    = ( l_44 [152] & !i[1704]) | ( l_44 [153] &  i[1704]);
assign l_43[78]    = ( l_44 [154] & !i[1704]) | ( l_44 [155] &  i[1704]);
assign l_43[79]    = ( l_44 [156] & !i[1704]) | ( l_44 [157] &  i[1704]);
assign l_43[80]    = ( l_44 [158] & !i[1704]) | ( l_44 [159] &  i[1704]);
assign l_43[81]    = ( l_44 [160] & !i[1704]) | ( l_44 [161] &  i[1704]);
assign l_43[82]    = ( l_44 [162] & !i[1704]) | ( l_44 [163] &  i[1704]);
assign l_43[83]    = ( l_44 [164] & !i[1704]) | ( l_44 [165] &  i[1704]);
assign l_43[84]    = ( l_44 [166] & !i[1704]) | ( l_44 [167] &  i[1704]);
assign l_43[85]    = ( l_44 [168] & !i[1704]) | ( l_44 [169] &  i[1704]);
assign l_43[86]    = ( l_44 [170] & !i[1704]) | ( l_44 [171] &  i[1704]);
assign l_43[87]    = ( l_44 [172] & !i[1704]) | ( l_44 [173] &  i[1704]);
assign l_43[88]    = ( l_44 [174] & !i[1704]) | ( l_44 [175] &  i[1704]);
assign l_43[89]    = ( l_44 [176] & !i[1704]) | ( l_44 [177] &  i[1704]);
assign l_43[90]    = ( l_44 [178] & !i[1704]) | ( l_44 [179] &  i[1704]);
assign l_43[91]    = ( l_44 [180] & !i[1704]) | ( l_44 [181] &  i[1704]);
assign l_43[92]    = ( l_44 [182] & !i[1704]) | ( l_44 [183] &  i[1704]);
assign l_43[93]    = ( l_44 [184] & !i[1704]) | ( l_44 [185] &  i[1704]);
assign l_43[94]    = ( l_44 [186] & !i[1704]) | ( l_44 [187] &  i[1704]);
assign l_43[95]    = ( l_44 [188] & !i[1704]) | ( l_44 [189] &  i[1704]);
assign l_43[96]    = ( l_44 [190] & !i[1704]) | ( l_44 [191] &  i[1704]);
assign l_43[97]    = ( l_44 [192] & !i[1704]) | ( l_44 [193] &  i[1704]);
assign l_43[98]    = ( l_44 [194] & !i[1704]) | ( l_44 [195] &  i[1704]);
assign l_43[99]    = ( l_44 [196] & !i[1704]) | ( l_44 [197] &  i[1704]);
assign l_43[100]    = ( l_44 [198] & !i[1704]) | ( l_44 [199] &  i[1704]);
assign l_43[101]    = ( l_44 [200] & !i[1704]) | ( l_44 [201] &  i[1704]);
assign l_43[102]    = ( l_44 [202] & !i[1704]) | ( l_44 [203] &  i[1704]);
assign l_43[103]    = ( l_44 [204] & !i[1704]) | ( l_44 [205] &  i[1704]);
assign l_43[104]    = ( l_44 [206] & !i[1704]) | ( l_44 [207] &  i[1704]);
assign l_43[105]    = ( l_44 [208] & !i[1704]) | ( l_44 [209] &  i[1704]);
assign l_43[106]    = ( l_44 [210] & !i[1704]) | ( l_44 [211] &  i[1704]);
assign l_43[107]    = ( l_44 [212] & !i[1704]) | ( l_44 [213] &  i[1704]);
assign l_43[108]    = ( l_44 [214] & !i[1704]) | ( l_44 [215] &  i[1704]);
assign l_43[109]    = ( l_44 [216] & !i[1704]) | ( l_44 [217] &  i[1704]);
assign l_43[110]    = ( l_44 [218] & !i[1704]) | ( l_44 [219] &  i[1704]);
assign l_43[111]    = ( l_44 [220] & !i[1704]) | ( l_44 [221] &  i[1704]);
assign l_43[112]    = ( l_44 [222] & !i[1704]) | ( l_44 [223] &  i[1704]);
assign l_43[113]    = ( l_44 [224] & !i[1704]) | ( l_44 [225] &  i[1704]);
assign l_43[114]    = ( l_44 [226] & !i[1704]) | ( l_44 [227] &  i[1704]);
assign l_43[115]    = ( l_44 [228] & !i[1704]) | ( l_44 [229] &  i[1704]);
assign l_43[116]    = ( l_44 [230] & !i[1704]) | ( l_44 [231] &  i[1704]);
assign l_43[117]    = ( l_44 [232] & !i[1704]) | ( l_44 [233] &  i[1704]);
assign l_43[118]    = ( l_44 [234] & !i[1704]) | ( l_44 [235] &  i[1704]);
assign l_43[119]    = ( l_44 [236] & !i[1704]) | ( l_44 [237] &  i[1704]);
assign l_43[120]    = ( l_44 [238] & !i[1704]) | ( l_44 [239] &  i[1704]);
assign l_43[121]    = ( l_44 [240] & !i[1704]) | ( l_44 [241] &  i[1704]);
assign l_43[122]    = ( l_44 [242] & !i[1704]) | ( l_44 [243] &  i[1704]);
assign l_43[123]    = ( l_44 [244] & !i[1704]) | ( l_44 [245] &  i[1704]);
assign l_43[124]    = ( l_44 [246] & !i[1704]) | ( l_44 [247] &  i[1704]);
assign l_43[125]    = ( l_44 [248] & !i[1704]) | ( l_44 [249] &  i[1704]);
assign l_43[126]    = ( l_44 [250] & !i[1704]) | ( l_44 [251] &  i[1704]);
assign l_43[127]    = ( l_44 [252] & !i[1704]) | ( l_44 [253] &  i[1704]);
assign l_43[128]    = ( l_44 [254] & !i[1704]) | ( l_44 [255] &  i[1704]);
assign l_43[129]    = ( l_44 [256] & !i[1704]) | ( l_44 [257] &  i[1704]);
assign l_43[130]    = ( l_44 [258] & !i[1704]) | ( l_44 [259] &  i[1704]);
assign l_43[131]    = ( l_44 [258] & !i[1704]) | ( l_44 [260] &  i[1704]);
assign l_43[132]    = ( l_44 [258] & !i[1704]) | ( l_44 [261] &  i[1704]);
assign l_43[133]    = ( l_44 [258] & !i[1704]) | ( l_44 [262] &  i[1704]);
assign l_43[134]    = ( l_44 [258] & !i[1704]) | ( l_44 [263] &  i[1704]);
assign l_43[135]    = ( l_44 [258] & !i[1704]) | ( l_44 [264] &  i[1704]);
assign l_43[136]    = ( l_44 [258] & !i[1704]) | ( l_44 [265] &  i[1704]);
assign l_43[137]    = ( l_44 [258] & !i[1704]) | ( l_44 [266] &  i[1704]);
assign l_43[138]    = ( l_44 [267] & !i[1704]);
assign l_43[139]    = ( l_44 [268] & !i[1704]);
assign l_43[140]    = ( l_44 [269] & !i[1704]);
assign l_43[141]    = ( l_44 [270] & !i[1704]);
assign l_43[142]    = ( l_44 [271] & !i[1704]);
assign l_43[143]    = ( l_44 [272] & !i[1704]);
assign l_43[144]    = ( l_44 [267] &  i[1704]);
assign l_43[145]    = ( l_44 [0] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[146]    = ( l_44 [267]);
assign l_43[147]    = ( l_44 [268] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[148]    = ( l_44 [269] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[149]    = ( l_44 [270] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[150]    = ( l_44 [271] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[151]    = ( l_44 [272] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[152]    = ( l_44 [0] &  i[1704]);
assign l_43[153]    = ( l_44 [0]);
assign l_43[154]    = ( l_44 [267] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[155]    = ( l_44 [268] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[156]    = ( l_44 [269] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[157]    = ( l_44 [270] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[158]    = ( l_44 [271] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[159]    = ( l_44 [272] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[160]    = ( l_44 [268] &  i[1704]);
assign l_43[161]    = ( l_44 [0] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[162]    = ( l_44 [267] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[163]    = ( l_44 [268]);
assign l_43[164]    = ( l_44 [269] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[165]    = ( l_44 [270] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[166]    = ( l_44 [271] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[167]    = ( l_44 [272] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[168]    = ( l_44 [273] &  i[1704]);
assign l_43[169]    = ( l_44 [0] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[170]    = ( l_44 [267] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[171]    = ( l_44 [268] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[172]    = ( l_44 [269] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[173]    = ( l_44 [270] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[174]    = ( l_44 [271] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[175]    = ( l_44 [272] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[176]    = ( l_44 [274] &  i[1704]);
assign l_43[177]    = ( l_44 [0] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[178]    = ( l_44 [267] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[179]    = ( l_44 [268] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[180]    = ( l_44 [269] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[181]    = ( l_44 [270] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[182]    = ( l_44 [271] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[183]    = ( l_44 [272] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[184]    = ( l_44 [275] &  i[1704]);
assign l_43[185]    = ( l_44 [0] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[186]    = ( l_44 [267] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[187]    = ( l_44 [268] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[188]    = ( l_44 [269] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[189]    = ( l_44 [270] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[190]    = ( l_44 [271] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[191]    = ( l_44 [272] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[192]    = ( l_44 [276] &  i[1704]);
assign l_43[193]    = ( l_44 [0] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[194]    = ( l_44 [267] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[195]    = ( l_44 [268] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[196]    = ( l_44 [269] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[197]    = ( l_44 [270] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[198]    = ( l_44 [271] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[199]    = ( l_44 [272] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[200]    = ( l_44 [269] &  i[1704]);
assign l_43[201]    = ( l_44 [0] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[202]    = ( l_44 [267] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[203]    = ( l_44 [268] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[204]    = ( l_44 [269]);
assign l_43[205]    = ( l_44 [270] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[206]    = ( l_44 [271] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[207]    = ( l_44 [272] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[208]    = ( l_44 [271] &  i[1704]);
assign l_43[209]    = ( l_44 [0] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[210]    = ( l_44 [267] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[211]    = ( l_44 [268] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[212]    = ( l_44 [269] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[213]    = ( l_44 [270] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[214]    = ( l_44 [271]);
assign l_43[215]    = ( l_44 [272] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[216]    = ( l_44 [270] &  i[1704]);
assign l_43[217]    = ( l_44 [0] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[218]    = ( l_44 [267] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[219]    = ( l_44 [268] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[220]    = ( l_44 [269] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[221]    = ( l_44 [270]);
assign l_43[222]    = ( l_44 [271] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[223]    = ( l_44 [272] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[224]    = ( l_44 [272] &  i[1704]);
assign l_43[225]    = ( l_44 [0] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[226]    = ( l_44 [267] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[227]    = ( l_44 [268] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[228]    = ( l_44 [269] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[229]    = ( l_44 [270] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[230]    = ( l_44 [271] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[231]    = ( l_44 [272]);
assign l_43[232]    = ( l_44 [277] &  i[1704]);
assign l_43[233]    = ( l_44 [0] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[234]    = ( l_44 [267] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[235]    = ( l_44 [268] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[236]    = ( l_44 [269] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[237]    = ( l_44 [270] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[238]    = ( l_44 [271] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[239]    = ( l_44 [272] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[240]    = ( l_44 [278] &  i[1704]);
assign l_43[241]    = ( l_44 [0] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[242]    = ( l_44 [267] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[243]    = ( l_44 [268] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[244]    = ( l_44 [269] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[245]    = ( l_44 [270] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[246]    = ( l_44 [271] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[247]    = ( l_44 [272] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[248]    = ( l_44 [279] &  i[1704]);
assign l_43[249]    = ( l_44 [0] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[250]    = ( l_44 [267] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[251]    = ( l_44 [268] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[252]    = ( l_44 [269] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[253]    = ( l_44 [270] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[254]    = ( l_44 [271] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[255]    = ( l_44 [272] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[256]    =  i[1704];
assign l_43[257]    = ( l_44 [0] & !i[1704]) | (      i[1704]);
assign l_43[258]    = ( l_44 [267] & !i[1704]) | (      i[1704]);
assign l_43[259]    = ( l_44 [268] & !i[1704]) | (      i[1704]);
assign l_43[260]    = ( l_44 [269] & !i[1704]) | (      i[1704]);
assign l_43[261]    = ( l_44 [270] & !i[1704]) | (      i[1704]);
assign l_43[262]    = ( l_44 [271] & !i[1704]) | (      i[1704]);
assign l_43[263]    = ( l_44 [272] & !i[1704]) | (      i[1704]);
assign l_43[264]    = ( l_44 [273] & !i[1704]);
assign l_43[265]    = ( l_44 [275] & !i[1704]);
assign l_43[266]    = ( l_44 [274] & !i[1704]);
assign l_43[267]    = ( l_44 [276] & !i[1704]);
assign l_43[268]    = ( l_44 [277] & !i[1704]);
assign l_43[269]    = ( l_44 [279] & !i[1704]);
assign l_43[270]    = ( l_44 [278] & !i[1704]);
assign l_43[271]    = !i[1704];
assign l_43[272]    = ( l_44 [273] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[273]    = ( l_44 [275] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[274]    = ( l_44 [274] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[275]    = ( l_44 [276] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[276]    = ( l_44 [277] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[277]    = ( l_44 [279] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[278]    = ( l_44 [278] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[279]    = (!i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[280]    = ( l_44 [273] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[281]    = ( l_44 [275] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[282]    = ( l_44 [274] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[283]    = ( l_44 [276] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[284]    = ( l_44 [277] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[285]    = ( l_44 [279] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[286]    = ( l_44 [278] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[287]    = (!i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[288]    = ( l_44 [273] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[289]    = ( l_44 [275] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[290]    = ( l_44 [274] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[291]    = ( l_44 [276] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[292]    = ( l_44 [277] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[293]    = ( l_44 [279] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[294]    = ( l_44 [278] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[295]    = (!i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[296]    = ( l_44 [273]);
assign l_43[297]    = ( l_44 [275] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[298]    = ( l_44 [274] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[299]    = ( l_44 [276] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[300]    = ( l_44 [277] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[301]    = ( l_44 [279] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[302]    = ( l_44 [278] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[303]    = (!i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[304]    = ( l_44 [273] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[305]    = ( l_44 [275] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[306]    = ( l_44 [274]);
assign l_43[307]    = ( l_44 [276] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[308]    = ( l_44 [277] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[309]    = ( l_44 [279] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[310]    = ( l_44 [278] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[311]    = (!i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[312]    = ( l_44 [273] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[313]    = ( l_44 [275]);
assign l_43[314]    = ( l_44 [274] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[315]    = ( l_44 [276] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[316]    = ( l_44 [277] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[317]    = ( l_44 [279] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[318]    = ( l_44 [278] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[319]    = (!i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[320]    = ( l_44 [273] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[321]    = ( l_44 [275] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[322]    = ( l_44 [274] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[323]    = ( l_44 [276]);
assign l_43[324]    = ( l_44 [277] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[325]    = ( l_44 [279] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[326]    = ( l_44 [278] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[327]    = (!i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[328]    = ( l_44 [273] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[329]    = ( l_44 [275] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[330]    = ( l_44 [274] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[331]    = ( l_44 [276] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[332]    = ( l_44 [277] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[333]    = ( l_44 [279] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[334]    = ( l_44 [278] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[335]    = (!i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[336]    = ( l_44 [273] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[337]    = ( l_44 [275] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[338]    = ( l_44 [274] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[339]    = ( l_44 [276] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[340]    = ( l_44 [277] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[341]    = ( l_44 [279] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[342]    = ( l_44 [278] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[343]    = (!i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[344]    = ( l_44 [273] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[345]    = ( l_44 [275] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[346]    = ( l_44 [274] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[347]    = ( l_44 [276] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[348]    = ( l_44 [277] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[349]    = ( l_44 [279] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[350]    = ( l_44 [278] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[351]    = (!i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[352]    = ( l_44 [273] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[353]    = ( l_44 [275] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[354]    = ( l_44 [274] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[355]    = ( l_44 [276] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[356]    = ( l_44 [277] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[357]    = ( l_44 [279] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[358]    = ( l_44 [278] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[359]    = (!i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[360]    = ( l_44 [273] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[361]    = ( l_44 [275] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[362]    = ( l_44 [274] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[363]    = ( l_44 [276] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[364]    = ( l_44 [277]);
assign l_43[365]    = ( l_44 [279] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[366]    = ( l_44 [278] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[367]    = (!i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[368]    = ( l_44 [273] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[369]    = ( l_44 [275] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[370]    = ( l_44 [274] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[371]    = ( l_44 [276] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[372]    = ( l_44 [277] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[373]    = ( l_44 [279] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[374]    = ( l_44 [278]);
assign l_43[375]    = (!i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[376]    = ( l_44 [273] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[377]    = ( l_44 [275] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[378]    = ( l_44 [274] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[379]    = ( l_44 [276] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[380]    = ( l_44 [277] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[381]    = ( l_44 [279]);
assign l_43[382]    = ( l_44 [278] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[383]    = (!i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[384]    = ( l_44 [273] & !i[1704]) | (      i[1704]);
assign l_43[385]    = ( l_44 [275] & !i[1704]) | (      i[1704]);
assign l_43[386]    = ( l_44 [274] & !i[1704]) | (      i[1704]);
assign l_43[387]    = ( l_44 [276] & !i[1704]) | (      i[1704]);
assign l_43[388]    = ( l_44 [277] & !i[1704]) | (      i[1704]);
assign l_43[389]    = ( l_44 [279] & !i[1704]) | (      i[1704]);
assign l_43[390]    = ( l_44 [278] & !i[1704]) | (      i[1704]);
assign l_43[391]    = ( l_44 [280] & !i[1704]) | ( l_44 [259] &  i[1704]);
assign l_43[392]    = ( l_44 [280] & !i[1704]) | ( l_44 [260] &  i[1704]);
assign l_43[393]    = ( l_44 [280] & !i[1704]) | ( l_44 [261] &  i[1704]);
assign l_43[394]    = ( l_44 [280] & !i[1704]) | ( l_44 [262] &  i[1704]);
assign l_43[395]    = ( l_44 [280] & !i[1704]) | ( l_44 [263] &  i[1704]);
assign l_43[396]    = ( l_44 [280] & !i[1704]) | ( l_44 [264] &  i[1704]);
assign l_43[397]    = ( l_44 [280] & !i[1704]) | ( l_44 [265] &  i[1704]);
assign l_43[398]    = ( l_44 [280] & !i[1704]) | ( l_44 [266] &  i[1704]);
assign l_43[399]    = ( l_44 [281] & !i[1704]);
assign l_43[400]    = ( l_44 [281] & !i[1704]) | ( l_44 [0] &  i[1704]);
assign l_43[401]    = ( l_44 [281] & !i[1704]) | ( l_44 [267] &  i[1704]);
assign l_43[402]    = ( l_44 [281] & !i[1704]) | ( l_44 [268] &  i[1704]);
assign l_43[403]    = ( l_44 [281] & !i[1704]) | ( l_44 [269] &  i[1704]);
assign l_43[404]    = ( l_44 [281] & !i[1704]) | ( l_44 [270] &  i[1704]);
assign l_43[405]    = ( l_44 [281] & !i[1704]) | ( l_44 [271] &  i[1704]);
assign l_43[406]    = ( l_44 [281] & !i[1704]) | ( l_44 [272] &  i[1704]);
assign l_43[407]    = ( l_44 [281] & !i[1704]) | ( l_44 [273] &  i[1704]);
assign l_43[408]    = ( l_44 [281] & !i[1704]) | ( l_44 [275] &  i[1704]);
assign l_43[409]    = ( l_44 [281] & !i[1704]) | ( l_44 [274] &  i[1704]);
assign l_43[410]    = ( l_44 [281] & !i[1704]) | ( l_44 [276] &  i[1704]);
assign l_43[411]    = ( l_44 [281] & !i[1704]) | ( l_44 [277] &  i[1704]);
assign l_43[412]    = ( l_44 [281] & !i[1704]) | ( l_44 [279] &  i[1704]);
assign l_43[413]    = ( l_44 [281] & !i[1704]) | ( l_44 [278] &  i[1704]);
assign l_43[414]    = ( l_44 [281] & !i[1704]) | (      i[1704]);
assign l_44[0]    = ( l_45 [0] & !i[1706]);
assign l_44[1]    = ( l_45 [1] & !i[1706]) | ( l_45 [2] &  i[1706]);
assign l_44[2]    = ( l_45 [3] & !i[1706]) | ( l_45 [4] &  i[1706]);
assign l_44[3]    = ( l_45 [5] & !i[1706]) | ( l_45 [6] &  i[1706]);
assign l_44[4]    = ( l_45 [7] & !i[1706]) | ( l_45 [8] &  i[1706]);
assign l_44[5]    = ( l_45 [9] & !i[1706]) | ( l_45 [10] &  i[1706]);
assign l_44[6]    = ( l_45 [11] & !i[1706]) | ( l_45 [12] &  i[1706]);
assign l_44[7]    = ( l_45 [13] & !i[1706]) | ( l_45 [14] &  i[1706]);
assign l_44[8]    = ( l_45 [15] & !i[1706]) | ( l_45 [16] &  i[1706]);
assign l_44[9]    = ( l_45 [17] & !i[1706]) | ( l_45 [18] &  i[1706]);
assign l_44[10]    = ( l_45 [19] & !i[1706]) | ( l_45 [20] &  i[1706]);
assign l_44[11]    = ( l_45 [21] & !i[1706]) | ( l_45 [22] &  i[1706]);
assign l_44[12]    = ( l_45 [23] & !i[1706]) | ( l_45 [24] &  i[1706]);
assign l_44[13]    = ( l_45 [25] & !i[1706]) | ( l_45 [26] &  i[1706]);
assign l_44[14]    = ( l_45 [27] & !i[1706]) | ( l_45 [28] &  i[1706]);
assign l_44[15]    = ( l_45 [29] & !i[1706]) | ( l_45 [30] &  i[1706]);
assign l_44[16]    = ( l_45 [31] & !i[1706]) | ( l_45 [32] &  i[1706]);
assign l_44[17]    = ( l_45 [33] & !i[1706]) | ( l_45 [34] &  i[1706]);
assign l_44[18]    = ( l_45 [35] & !i[1706]) | ( l_45 [36] &  i[1706]);
assign l_44[19]    = ( l_45 [37] & !i[1706]) | ( l_45 [38] &  i[1706]);
assign l_44[20]    = ( l_45 [39] & !i[1706]) | ( l_45 [40] &  i[1706]);
assign l_44[21]    = ( l_45 [41] & !i[1706]) | ( l_45 [42] &  i[1706]);
assign l_44[22]    = ( l_45 [43] & !i[1706]) | ( l_45 [44] &  i[1706]);
assign l_44[23]    = ( l_45 [45] & !i[1706]) | ( l_45 [46] &  i[1706]);
assign l_44[24]    = ( l_45 [47] & !i[1706]) | ( l_45 [48] &  i[1706]);
assign l_44[25]    = ( l_45 [49] & !i[1706]) | ( l_45 [50] &  i[1706]);
assign l_44[26]    = ( l_45 [51] & !i[1706]) | ( l_45 [52] &  i[1706]);
assign l_44[27]    = ( l_45 [53] & !i[1706]) | ( l_45 [54] &  i[1706]);
assign l_44[28]    = ( l_45 [55] & !i[1706]) | ( l_45 [56] &  i[1706]);
assign l_44[29]    = ( l_45 [57] & !i[1706]) | ( l_45 [58] &  i[1706]);
assign l_44[30]    = ( l_45 [59] & !i[1706]) | ( l_45 [60] &  i[1706]);
assign l_44[31]    = ( l_45 [61] & !i[1706]) | ( l_45 [62] &  i[1706]);
assign l_44[32]    = ( l_45 [63] & !i[1706]) | ( l_45 [64] &  i[1706]);
assign l_44[33]    = ( l_45 [65] & !i[1706]) | ( l_45 [66] &  i[1706]);
assign l_44[34]    = ( l_45 [67] & !i[1706]) | ( l_45 [68] &  i[1706]);
assign l_44[35]    = ( l_45 [69] & !i[1706]) | ( l_45 [70] &  i[1706]);
assign l_44[36]    = ( l_45 [71] & !i[1706]) | ( l_45 [72] &  i[1706]);
assign l_44[37]    = ( l_45 [73] & !i[1706]) | ( l_45 [74] &  i[1706]);
assign l_44[38]    = ( l_45 [75] & !i[1706]) | ( l_45 [76] &  i[1706]);
assign l_44[39]    = ( l_45 [77] & !i[1706]) | ( l_45 [78] &  i[1706]);
assign l_44[40]    = ( l_45 [79] & !i[1706]) | ( l_45 [80] &  i[1706]);
assign l_44[41]    = ( l_45 [81] & !i[1706]) | ( l_45 [82] &  i[1706]);
assign l_44[42]    = ( l_45 [83] & !i[1706]) | ( l_45 [84] &  i[1706]);
assign l_44[43]    = ( l_45 [85] & !i[1706]) | ( l_45 [86] &  i[1706]);
assign l_44[44]    = ( l_45 [87] & !i[1706]) | ( l_45 [88] &  i[1706]);
assign l_44[45]    = ( l_45 [89] & !i[1706]) | ( l_45 [90] &  i[1706]);
assign l_44[46]    = ( l_45 [91] & !i[1706]) | ( l_45 [92] &  i[1706]);
assign l_44[47]    = ( l_45 [93] & !i[1706]) | ( l_45 [94] &  i[1706]);
assign l_44[48]    = ( l_45 [95] & !i[1706]) | ( l_45 [96] &  i[1706]);
assign l_44[49]    = ( l_45 [97] & !i[1706]) | ( l_45 [98] &  i[1706]);
assign l_44[50]    = ( l_45 [99] & !i[1706]) | ( l_45 [100] &  i[1706]);
assign l_44[51]    = ( l_45 [101] & !i[1706]) | ( l_45 [102] &  i[1706]);
assign l_44[52]    = ( l_45 [103] & !i[1706]) | ( l_45 [104] &  i[1706]);
assign l_44[53]    = ( l_45 [105] & !i[1706]) | ( l_45 [106] &  i[1706]);
assign l_44[54]    = ( l_45 [107] & !i[1706]) | ( l_45 [108] &  i[1706]);
assign l_44[55]    = ( l_45 [109] & !i[1706]) | ( l_45 [110] &  i[1706]);
assign l_44[56]    = ( l_45 [111] & !i[1706]) | ( l_45 [112] &  i[1706]);
assign l_44[57]    = ( l_45 [113] & !i[1706]) | ( l_45 [114] &  i[1706]);
assign l_44[58]    = ( l_45 [115] & !i[1706]) | ( l_45 [116] &  i[1706]);
assign l_44[59]    = ( l_45 [117] & !i[1706]) | ( l_45 [118] &  i[1706]);
assign l_44[60]    = ( l_45 [119] & !i[1706]) | ( l_45 [120] &  i[1706]);
assign l_44[61]    = ( l_45 [121] & !i[1706]) | ( l_45 [122] &  i[1706]);
assign l_44[62]    = ( l_45 [123] & !i[1706]) | ( l_45 [124] &  i[1706]);
assign l_44[63]    = ( l_45 [125] & !i[1706]) | ( l_45 [126] &  i[1706]);
assign l_44[64]    = ( l_45 [127] & !i[1706]) | ( l_45 [128] &  i[1706]);
assign l_44[65]    = ( l_45 [2] & !i[1706]) | ( l_45 [129] &  i[1706]);
assign l_44[66]    = ( l_45 [4] & !i[1706]) | ( l_45 [130] &  i[1706]);
assign l_44[67]    = ( l_45 [6] & !i[1706]) | ( l_45 [131] &  i[1706]);
assign l_44[68]    = ( l_45 [8] & !i[1706]) | ( l_45 [132] &  i[1706]);
assign l_44[69]    = ( l_45 [10] & !i[1706]) | ( l_45 [133] &  i[1706]);
assign l_44[70]    = ( l_45 [12] & !i[1706]) | ( l_45 [134] &  i[1706]);
assign l_44[71]    = ( l_45 [14] & !i[1706]) | ( l_45 [135] &  i[1706]);
assign l_44[72]    = ( l_45 [16] & !i[1706]) | ( l_45 [136] &  i[1706]);
assign l_44[73]    = ( l_45 [18] & !i[1706]) | ( l_45 [137] &  i[1706]);
assign l_44[74]    = ( l_45 [20] & !i[1706]) | ( l_45 [138] &  i[1706]);
assign l_44[75]    = ( l_45 [22] & !i[1706]) | ( l_45 [139] &  i[1706]);
assign l_44[76]    = ( l_45 [24] & !i[1706]) | ( l_45 [140] &  i[1706]);
assign l_44[77]    = ( l_45 [26] & !i[1706]) | ( l_45 [141] &  i[1706]);
assign l_44[78]    = ( l_45 [28] & !i[1706]) | ( l_45 [142] &  i[1706]);
assign l_44[79]    = ( l_45 [30] & !i[1706]) | ( l_45 [143] &  i[1706]);
assign l_44[80]    = ( l_45 [32] & !i[1706]) | ( l_45 [144] &  i[1706]);
assign l_44[81]    = ( l_45 [34] & !i[1706]) | ( l_45 [145] &  i[1706]);
assign l_44[82]    = ( l_45 [36] & !i[1706]) | ( l_45 [146] &  i[1706]);
assign l_44[83]    = ( l_45 [38] & !i[1706]) | ( l_45 [147] &  i[1706]);
assign l_44[84]    = ( l_45 [40] & !i[1706]) | ( l_45 [148] &  i[1706]);
assign l_44[85]    = ( l_45 [42] & !i[1706]) | ( l_45 [149] &  i[1706]);
assign l_44[86]    = ( l_45 [44] & !i[1706]) | ( l_45 [150] &  i[1706]);
assign l_44[87]    = ( l_45 [46] & !i[1706]) | ( l_45 [151] &  i[1706]);
assign l_44[88]    = ( l_45 [48] & !i[1706]) | ( l_45 [152] &  i[1706]);
assign l_44[89]    = ( l_45 [50] & !i[1706]) | ( l_45 [153] &  i[1706]);
assign l_44[90]    = ( l_45 [52] & !i[1706]) | ( l_45 [154] &  i[1706]);
assign l_44[91]    = ( l_45 [54] & !i[1706]) | ( l_45 [155] &  i[1706]);
assign l_44[92]    = ( l_45 [56] & !i[1706]) | ( l_45 [156] &  i[1706]);
assign l_44[93]    = ( l_45 [58] & !i[1706]) | ( l_45 [157] &  i[1706]);
assign l_44[94]    = ( l_45 [60] & !i[1706]) | ( l_45 [158] &  i[1706]);
assign l_44[95]    = ( l_45 [62] & !i[1706]) | ( l_45 [159] &  i[1706]);
assign l_44[96]    = ( l_45 [64] & !i[1706]) | ( l_45 [160] &  i[1706]);
assign l_44[97]    = ( l_45 [66] & !i[1706]) | ( l_45 [161] &  i[1706]);
assign l_44[98]    = ( l_45 [68] & !i[1706]) | ( l_45 [162] &  i[1706]);
assign l_44[99]    = ( l_45 [70] & !i[1706]) | ( l_45 [163] &  i[1706]);
assign l_44[100]    = ( l_45 [72] & !i[1706]) | ( l_45 [164] &  i[1706]);
assign l_44[101]    = ( l_45 [74] & !i[1706]) | ( l_45 [165] &  i[1706]);
assign l_44[102]    = ( l_45 [76] & !i[1706]) | ( l_45 [166] &  i[1706]);
assign l_44[103]    = ( l_45 [78] & !i[1706]) | ( l_45 [167] &  i[1706]);
assign l_44[104]    = ( l_45 [80] & !i[1706]) | ( l_45 [168] &  i[1706]);
assign l_44[105]    = ( l_45 [82] & !i[1706]) | ( l_45 [169] &  i[1706]);
assign l_44[106]    = ( l_45 [84] & !i[1706]) | ( l_45 [170] &  i[1706]);
assign l_44[107]    = ( l_45 [86] & !i[1706]) | ( l_45 [171] &  i[1706]);
assign l_44[108]    = ( l_45 [88] & !i[1706]) | ( l_45 [172] &  i[1706]);
assign l_44[109]    = ( l_45 [90] & !i[1706]) | ( l_45 [173] &  i[1706]);
assign l_44[110]    = ( l_45 [92] & !i[1706]) | ( l_45 [174] &  i[1706]);
assign l_44[111]    = ( l_45 [94] & !i[1706]) | ( l_45 [175] &  i[1706]);
assign l_44[112]    = ( l_45 [96] & !i[1706]) | ( l_45 [176] &  i[1706]);
assign l_44[113]    = ( l_45 [98] & !i[1706]) | ( l_45 [177] &  i[1706]);
assign l_44[114]    = ( l_45 [100] & !i[1706]) | ( l_45 [178] &  i[1706]);
assign l_44[115]    = ( l_45 [102] & !i[1706]) | ( l_45 [179] &  i[1706]);
assign l_44[116]    = ( l_45 [104] & !i[1706]) | ( l_45 [180] &  i[1706]);
assign l_44[117]    = ( l_45 [106] & !i[1706]) | ( l_45 [181] &  i[1706]);
assign l_44[118]    = ( l_45 [108] & !i[1706]) | ( l_45 [182] &  i[1706]);
assign l_44[119]    = ( l_45 [110] & !i[1706]) | ( l_45 [183] &  i[1706]);
assign l_44[120]    = ( l_45 [112] & !i[1706]) | ( l_45 [184] &  i[1706]);
assign l_44[121]    = ( l_45 [114] & !i[1706]) | ( l_45 [185] &  i[1706]);
assign l_44[122]    = ( l_45 [116] & !i[1706]) | ( l_45 [186] &  i[1706]);
assign l_44[123]    = ( l_45 [118] & !i[1706]) | ( l_45 [187] &  i[1706]);
assign l_44[124]    = ( l_45 [120] & !i[1706]) | ( l_45 [188] &  i[1706]);
assign l_44[125]    = ( l_45 [122] & !i[1706]) | ( l_45 [189] &  i[1706]);
assign l_44[126]    = ( l_45 [124] & !i[1706]) | ( l_45 [190] &  i[1706]);
assign l_44[127]    = ( l_45 [126] & !i[1706]) | ( l_45 [191] &  i[1706]);
assign l_44[128]    = ( l_45 [128] & !i[1706]) | ( l_45 [192] &  i[1706]);
assign l_44[129]    = ( l_45 [193] & !i[1706]) | ( l_45 [194] &  i[1706]);
assign l_44[130]    = ( l_45 [195] & !i[1706]) | ( l_45 [196] &  i[1706]);
assign l_44[131]    = ( l_45 [197] & !i[1706]) | ( l_45 [198] &  i[1706]);
assign l_44[132]    = ( l_45 [199] & !i[1706]) | ( l_45 [200] &  i[1706]);
assign l_44[133]    = ( l_45 [201] & !i[1706]) | ( l_45 [202] &  i[1706]);
assign l_44[134]    = ( l_45 [203] & !i[1706]) | ( l_45 [204] &  i[1706]);
assign l_44[135]    = ( l_45 [205] & !i[1706]) | ( l_45 [206] &  i[1706]);
assign l_44[136]    = ( l_45 [207] & !i[1706]) | ( l_45 [208] &  i[1706]);
assign l_44[137]    = ( l_45 [209] & !i[1706]) | ( l_45 [210] &  i[1706]);
assign l_44[138]    = ( l_45 [211] & !i[1706]) | ( l_45 [212] &  i[1706]);
assign l_44[139]    = ( l_45 [213] & !i[1706]) | ( l_45 [214] &  i[1706]);
assign l_44[140]    = ( l_45 [215] & !i[1706]) | ( l_45 [216] &  i[1706]);
assign l_44[141]    = ( l_45 [217] & !i[1706]) | ( l_45 [218] &  i[1706]);
assign l_44[142]    = ( l_45 [219] & !i[1706]) | ( l_45 [220] &  i[1706]);
assign l_44[143]    = ( l_45 [221] & !i[1706]) | ( l_45 [222] &  i[1706]);
assign l_44[144]    = ( l_45 [223] & !i[1706]) | ( l_45 [224] &  i[1706]);
assign l_44[145]    = ( l_45 [225]);
assign l_44[146]    = ( l_45 [226] & !i[1706]) | ( l_45 [227] &  i[1706]);
assign l_44[147]    = ( l_45 [228] & !i[1706]) | ( l_45 [229] &  i[1706]);
assign l_44[148]    = ( l_45 [230] & !i[1706]) | ( l_45 [231] &  i[1706]);
assign l_44[149]    = ( l_45 [232] & !i[1706]) | ( l_45 [233] &  i[1706]);
assign l_44[150]    = ( l_45 [234] & !i[1706]) | ( l_45 [235] &  i[1706]);
assign l_44[151]    = ( l_45 [236] & !i[1706]) | ( l_45 [237] &  i[1706]);
assign l_44[152]    = ( l_45 [238] & !i[1706]) | ( l_45 [239] &  i[1706]);
assign l_44[153]    = ( l_45 [240] & !i[1706]) | ( l_45 [241] &  i[1706]);
assign l_44[154]    = ( l_45 [242] & !i[1706]) | ( l_45 [243] &  i[1706]);
assign l_44[155]    = ( l_45 [244] & !i[1706]) | ( l_45 [245] &  i[1706]);
assign l_44[156]    = ( l_45 [246] & !i[1706]) | ( l_45 [247] &  i[1706]);
assign l_44[157]    = ( l_45 [248] & !i[1706]) | ( l_45 [249] &  i[1706]);
assign l_44[158]    = ( l_45 [250] & !i[1706]) | ( l_45 [251] &  i[1706]);
assign l_44[159]    = ( l_45 [252] & !i[1706]) | ( l_45 [253] &  i[1706]);
assign l_44[160]    = ( l_45 [254] & !i[1706]) | ( l_45 [255] &  i[1706]);
assign l_44[161]    = ( l_45 [256] & !i[1706]) | ( l_45 [257] &  i[1706]);
assign l_44[162]    = ( l_45 [258] & !i[1706]) | ( l_45 [259] &  i[1706]);
assign l_44[163]    = ( l_45 [260] & !i[1706]) | ( l_45 [261] &  i[1706]);
assign l_44[164]    = ( l_45 [262] & !i[1706]) | ( l_45 [263] &  i[1706]);
assign l_44[165]    = ( l_45 [264] & !i[1706]) | ( l_45 [265] &  i[1706]);
assign l_44[166]    = ( l_45 [266] & !i[1706]) | ( l_45 [267] &  i[1706]);
assign l_44[167]    = ( l_45 [268] & !i[1706]) | ( l_45 [269] &  i[1706]);
assign l_44[168]    = ( l_45 [270] & !i[1706]) | ( l_45 [271] &  i[1706]);
assign l_44[169]    = ( l_45 [272] & !i[1706]) | ( l_45 [273] &  i[1706]);
assign l_44[170]    = ( l_45 [274] & !i[1706]) | ( l_45 [275] &  i[1706]);
assign l_44[171]    = ( l_45 [276] & !i[1706]) | ( l_45 [277] &  i[1706]);
assign l_44[172]    = ( l_45 [278] & !i[1706]) | ( l_45 [279] &  i[1706]);
assign l_44[173]    = ( l_45 [280] & !i[1706]) | ( l_45 [281] &  i[1706]);
assign l_44[174]    = ( l_45 [282] & !i[1706]) | ( l_45 [283] &  i[1706]);
assign l_44[175]    = ( l_45 [284] & !i[1706]) | ( l_45 [285] &  i[1706]);
assign l_44[176]    = ( l_45 [286] & !i[1706]) | ( l_45 [287] &  i[1706]);
assign l_44[177]    = ( l_45 [288] & !i[1706]) | ( l_45 [289] &  i[1706]);
assign l_44[178]    = ( l_45 [290] & !i[1706]) | ( l_45 [291] &  i[1706]);
assign l_44[179]    = ( l_45 [292] & !i[1706]) | ( l_45 [293] &  i[1706]);
assign l_44[180]    = ( l_45 [294] & !i[1706]) | ( l_45 [295] &  i[1706]);
assign l_44[181]    = ( l_45 [296] & !i[1706]) | ( l_45 [297] &  i[1706]);
assign l_44[182]    = ( l_45 [298] & !i[1706]) | ( l_45 [299] &  i[1706]);
assign l_44[183]    = ( l_45 [300] & !i[1706]) | ( l_45 [301] &  i[1706]);
assign l_44[184]    = ( l_45 [302] & !i[1706]) | ( l_45 [303] &  i[1706]);
assign l_44[185]    = ( l_45 [304] & !i[1706]) | ( l_45 [305] &  i[1706]);
assign l_44[186]    = ( l_45 [306] & !i[1706]) | ( l_45 [307] &  i[1706]);
assign l_44[187]    = ( l_45 [308] & !i[1706]) | ( l_45 [309] &  i[1706]);
assign l_44[188]    = ( l_45 [310] & !i[1706]) | ( l_45 [311] &  i[1706]);
assign l_44[189]    = ( l_45 [312] & !i[1706]) | ( l_45 [313] &  i[1706]);
assign l_44[190]    = ( l_45 [314] & !i[1706]) | ( l_45 [315] &  i[1706]);
assign l_44[191]    = ( l_45 [316] & !i[1706]) | ( l_45 [317] &  i[1706]);
assign l_44[192]    = ( l_45 [318] & !i[1706]) | ( l_45 [319] &  i[1706]);
assign l_44[193]    = ( l_45 [320] & !i[1706]) | ( l_45 [321] &  i[1706]);
assign l_44[194]    = ( l_45 [194] & !i[1706]) | ( l_45 [322] &  i[1706]);
assign l_44[195]    = ( l_45 [196] & !i[1706]) | ( l_45 [323] &  i[1706]);
assign l_44[196]    = ( l_45 [198] & !i[1706]) | ( l_45 [324] &  i[1706]);
assign l_44[197]    = ( l_45 [200] & !i[1706]) | ( l_45 [325] &  i[1706]);
assign l_44[198]    = ( l_45 [202] & !i[1706]) | ( l_45 [326] &  i[1706]);
assign l_44[199]    = ( l_45 [204] & !i[1706]) | ( l_45 [327] &  i[1706]);
assign l_44[200]    = ( l_45 [206] & !i[1706]) | ( l_45 [328] &  i[1706]);
assign l_44[201]    = ( l_45 [208] & !i[1706]) | ( l_45 [329] &  i[1706]);
assign l_44[202]    = ( l_45 [210] & !i[1706]) | ( l_45 [330] &  i[1706]);
assign l_44[203]    = ( l_45 [212] & !i[1706]) | ( l_45 [331] &  i[1706]);
assign l_44[204]    = ( l_45 [214] & !i[1706]) | ( l_45 [332] &  i[1706]);
assign l_44[205]    = ( l_45 [216] & !i[1706]) | ( l_45 [333] &  i[1706]);
assign l_44[206]    = ( l_45 [218] & !i[1706]) | ( l_45 [334] &  i[1706]);
assign l_44[207]    = ( l_45 [220] & !i[1706]) | ( l_45 [335] &  i[1706]);
assign l_44[208]    = ( l_45 [222] & !i[1706]) | ( l_45 [336] &  i[1706]);
assign l_44[209]    = ( l_45 [224] & !i[1706]) | ( l_45 [337] &  i[1706]);
assign l_44[210]    = ( l_45 [227] & !i[1706]) | ( l_45 [338] &  i[1706]);
assign l_44[211]    = ( l_45 [229] & !i[1706]) | ( l_45 [339] &  i[1706]);
assign l_44[212]    = ( l_45 [231] & !i[1706]) | ( l_45 [340] &  i[1706]);
assign l_44[213]    = ( l_45 [233] & !i[1706]) | ( l_45 [341] &  i[1706]);
assign l_44[214]    = ( l_45 [235] & !i[1706]) | ( l_45 [342] &  i[1706]);
assign l_44[215]    = ( l_45 [237] & !i[1706]) | ( l_45 [343] &  i[1706]);
assign l_44[216]    = ( l_45 [239] & !i[1706]) | ( l_45 [344] &  i[1706]);
assign l_44[217]    = ( l_45 [241] & !i[1706]) | ( l_45 [345] &  i[1706]);
assign l_44[218]    = ( l_45 [243] & !i[1706]) | ( l_45 [346] &  i[1706]);
assign l_44[219]    = ( l_45 [245] & !i[1706]) | ( l_45 [347] &  i[1706]);
assign l_44[220]    = ( l_45 [247] & !i[1706]) | ( l_45 [348] &  i[1706]);
assign l_44[221]    = ( l_45 [249] & !i[1706]) | ( l_45 [349] &  i[1706]);
assign l_44[222]    = ( l_45 [251] & !i[1706]) | ( l_45 [350] &  i[1706]);
assign l_44[223]    = ( l_45 [253] & !i[1706]) | ( l_45 [351] &  i[1706]);
assign l_44[224]    = ( l_45 [255] & !i[1706]) | ( l_45 [352] &  i[1706]);
assign l_44[225]    = ( l_45 [257] & !i[1706]) | ( l_45 [353] &  i[1706]);
assign l_44[226]    = ( l_45 [259] & !i[1706]) | ( l_45 [354] &  i[1706]);
assign l_44[227]    = ( l_45 [261] & !i[1706]) | ( l_45 [355] &  i[1706]);
assign l_44[228]    = ( l_45 [263] & !i[1706]) | ( l_45 [356] &  i[1706]);
assign l_44[229]    = ( l_45 [265] & !i[1706]) | ( l_45 [357] &  i[1706]);
assign l_44[230]    = ( l_45 [267] & !i[1706]) | ( l_45 [358] &  i[1706]);
assign l_44[231]    = ( l_45 [269] & !i[1706]) | ( l_45 [359] &  i[1706]);
assign l_44[232]    = ( l_45 [271] & !i[1706]) | ( l_45 [360] &  i[1706]);
assign l_44[233]    = ( l_45 [273] & !i[1706]) | ( l_45 [361] &  i[1706]);
assign l_44[234]    = ( l_45 [275] & !i[1706]) | ( l_45 [362] &  i[1706]);
assign l_44[235]    = ( l_45 [277] & !i[1706]) | ( l_45 [363] &  i[1706]);
assign l_44[236]    = ( l_45 [279] & !i[1706]) | ( l_45 [364] &  i[1706]);
assign l_44[237]    = ( l_45 [281] & !i[1706]) | ( l_45 [365] &  i[1706]);
assign l_44[238]    = ( l_45 [283] & !i[1706]) | ( l_45 [366] &  i[1706]);
assign l_44[239]    = ( l_45 [285] & !i[1706]) | ( l_45 [367] &  i[1706]);
assign l_44[240]    = ( l_45 [287] & !i[1706]) | ( l_45 [368] &  i[1706]);
assign l_44[241]    = ( l_45 [289] & !i[1706]) | ( l_45 [369] &  i[1706]);
assign l_44[242]    = ( l_45 [291] & !i[1706]) | ( l_45 [370] &  i[1706]);
assign l_44[243]    = ( l_45 [293] & !i[1706]) | ( l_45 [371] &  i[1706]);
assign l_44[244]    = ( l_45 [295] & !i[1706]) | ( l_45 [372] &  i[1706]);
assign l_44[245]    = ( l_45 [297] & !i[1706]) | ( l_45 [373] &  i[1706]);
assign l_44[246]    = ( l_45 [299] & !i[1706]) | ( l_45 [374] &  i[1706]);
assign l_44[247]    = ( l_45 [301] & !i[1706]) | ( l_45 [375] &  i[1706]);
assign l_44[248]    = ( l_45 [303] & !i[1706]) | ( l_45 [376] &  i[1706]);
assign l_44[249]    = ( l_45 [305] & !i[1706]) | ( l_45 [377] &  i[1706]);
assign l_44[250]    = ( l_45 [307] & !i[1706]) | ( l_45 [378] &  i[1706]);
assign l_44[251]    = ( l_45 [309] & !i[1706]) | ( l_45 [379] &  i[1706]);
assign l_44[252]    = ( l_45 [311] & !i[1706]) | ( l_45 [380] &  i[1706]);
assign l_44[253]    = ( l_45 [313] & !i[1706]) | ( l_45 [381] &  i[1706]);
assign l_44[254]    = ( l_45 [315] & !i[1706]) | ( l_45 [382] &  i[1706]);
assign l_44[255]    = ( l_45 [317] & !i[1706]) | ( l_45 [383] &  i[1706]);
assign l_44[256]    = ( l_45 [319] & !i[1706]) | ( l_45 [384] &  i[1706]);
assign l_44[257]    = ( l_45 [321] & !i[1706]) | ( l_45 [385] &  i[1706]);
assign l_44[258]    = ( l_45 [386] & !i[1706]) | ( l_45 [387] &  i[1706]);
assign l_44[259]    = ( l_45 [388] & !i[1706]);
assign l_44[260]    = ( l_45 [388] & !i[1706]) | ( l_45 [0] &  i[1706]);
assign l_44[261]    = ( l_45 [389] & !i[1706]);
assign l_44[262]    = ( l_45 [389] & !i[1706]) | ( l_45 [0] &  i[1706]);
assign l_44[263]    = ( l_45 [388] & !i[1706]) | ( l_45 [390] &  i[1706]);
assign l_44[264]    = ( l_45 [388] & !i[1706]) | (      i[1706]);
assign l_44[265]    = ( l_45 [389] & !i[1706]) | ( l_45 [390] &  i[1706]);
assign l_44[266]    = ( l_45 [389] & !i[1706]) | (      i[1706]);
assign l_44[267]    = ( l_45 [390] &  i[1706]);
assign l_44[268]    = ( l_45 [0] & !i[1706]) | ( l_45 [390] &  i[1706]);
assign l_44[269]    = ( l_45 [0] &  i[1706]);
assign l_44[270]    = ( l_45 [0]);
assign l_44[271]    =  i[1706];
assign l_44[272]    = ( l_45 [0] & !i[1706]) | (      i[1706]);
assign l_44[273]    = ( l_45 [390] & !i[1706]);
assign l_44[274]    = ( l_45 [390]);
assign l_44[275]    = !i[1706];
assign l_44[276]    = (!i[1706]) | ( l_45 [390] &  i[1706]);
assign l_44[277]    = ( l_45 [390] & !i[1706]) | ( l_45 [0] &  i[1706]);
assign l_44[278]    = ( l_45 [390] & !i[1706]) | (      i[1706]);
assign l_44[279]    = (!i[1706]) | ( l_45 [0] &  i[1706]);
assign l_44[280]    = ( l_45 [391] & !i[1706]) | ( l_45 [387] &  i[1706]);
assign l_44[281]    = ( l_45 [392] & !i[1706]) | ( l_45 [393] &  i[1706]);
assign l_45[0]    = !i[1705];
assign l_45[1]    = ( l_46 [0] & !i[1705]) | ( l_46 [1] &  i[1705]);
assign l_45[2]    = ( l_46 [2] & !i[1705]) | ( l_46 [3] &  i[1705]);
assign l_45[3]    = ( l_46 [4] & !i[1705]) | ( l_46 [5] &  i[1705]);
assign l_45[4]    = ( l_46 [6] & !i[1705]) | ( l_46 [7] &  i[1705]);
assign l_45[5]    = ( l_46 [8] & !i[1705]) | ( l_46 [9] &  i[1705]);
assign l_45[6]    = ( l_46 [10] & !i[1705]) | ( l_46 [11] &  i[1705]);
assign l_45[7]    = ( l_46 [12] & !i[1705]) | ( l_46 [13] &  i[1705]);
assign l_45[8]    = ( l_46 [14] & !i[1705]) | ( l_46 [15] &  i[1705]);
assign l_45[9]    = ( l_46 [16] & !i[1705]) | ( l_46 [17] &  i[1705]);
assign l_45[10]    = ( l_46 [18] & !i[1705]) | ( l_46 [19] &  i[1705]);
assign l_45[11]    = ( l_46 [20] & !i[1705]) | ( l_46 [21] &  i[1705]);
assign l_45[12]    = ( l_46 [22] & !i[1705]) | ( l_46 [23] &  i[1705]);
assign l_45[13]    = ( l_46 [24] & !i[1705]) | ( l_46 [25] &  i[1705]);
assign l_45[14]    = ( l_46 [26] & !i[1705]) | ( l_46 [27] &  i[1705]);
assign l_45[15]    = ( l_46 [28] & !i[1705]) | ( l_46 [29] &  i[1705]);
assign l_45[16]    = ( l_46 [30] & !i[1705]) | ( l_46 [31] &  i[1705]);
assign l_45[17]    = ( l_46 [32] & !i[1705]) | ( l_46 [33] &  i[1705]);
assign l_45[18]    = ( l_46 [34] & !i[1705]) | ( l_46 [35] &  i[1705]);
assign l_45[19]    = ( l_46 [36] & !i[1705]) | ( l_46 [37] &  i[1705]);
assign l_45[20]    = ( l_46 [38] & !i[1705]) | ( l_46 [39] &  i[1705]);
assign l_45[21]    = ( l_46 [40] & !i[1705]) | ( l_46 [41] &  i[1705]);
assign l_45[22]    = ( l_46 [42] & !i[1705]) | ( l_46 [43] &  i[1705]);
assign l_45[23]    = ( l_46 [44] & !i[1705]) | ( l_46 [45] &  i[1705]);
assign l_45[24]    = ( l_46 [46] & !i[1705]) | ( l_46 [47] &  i[1705]);
assign l_45[25]    = ( l_46 [48] & !i[1705]) | ( l_46 [49] &  i[1705]);
assign l_45[26]    = ( l_46 [50] & !i[1705]) | ( l_46 [51] &  i[1705]);
assign l_45[27]    = ( l_46 [52] & !i[1705]) | ( l_46 [53] &  i[1705]);
assign l_45[28]    = ( l_46 [54] & !i[1705]) | ( l_46 [55] &  i[1705]);
assign l_45[29]    = ( l_46 [56] & !i[1705]) | ( l_46 [57] &  i[1705]);
assign l_45[30]    = ( l_46 [58] & !i[1705]) | ( l_46 [59] &  i[1705]);
assign l_45[31]    = ( l_46 [60] & !i[1705]) | ( l_46 [61] &  i[1705]);
assign l_45[32]    = ( l_46 [62] & !i[1705]) | ( l_46 [63] &  i[1705]);
assign l_45[33]    = ( l_46 [64] & !i[1705]) | ( l_46 [65] &  i[1705]);
assign l_45[34]    = ( l_46 [66] & !i[1705]) | ( l_46 [67] &  i[1705]);
assign l_45[35]    = ( l_46 [68] & !i[1705]) | ( l_46 [69] &  i[1705]);
assign l_45[36]    = ( l_46 [70] & !i[1705]) | ( l_46 [71] &  i[1705]);
assign l_45[37]    = ( l_46 [72] & !i[1705]) | ( l_46 [73] &  i[1705]);
assign l_45[38]    = ( l_46 [74] & !i[1705]) | ( l_46 [75] &  i[1705]);
assign l_45[39]    = ( l_46 [76] & !i[1705]) | ( l_46 [77] &  i[1705]);
assign l_45[40]    = ( l_46 [78] & !i[1705]) | ( l_46 [79] &  i[1705]);
assign l_45[41]    = ( l_46 [80] & !i[1705]) | ( l_46 [81] &  i[1705]);
assign l_45[42]    = ( l_46 [82] & !i[1705]) | ( l_46 [83] &  i[1705]);
assign l_45[43]    = ( l_46 [84] & !i[1705]) | ( l_46 [85] &  i[1705]);
assign l_45[44]    = ( l_46 [86] & !i[1705]) | ( l_46 [87] &  i[1705]);
assign l_45[45]    = ( l_46 [88] & !i[1705]) | ( l_46 [89] &  i[1705]);
assign l_45[46]    = ( l_46 [90] & !i[1705]) | ( l_46 [91] &  i[1705]);
assign l_45[47]    = ( l_46 [92] & !i[1705]) | ( l_46 [93] &  i[1705]);
assign l_45[48]    = ( l_46 [94] & !i[1705]) | ( l_46 [95] &  i[1705]);
assign l_45[49]    = ( l_46 [96] & !i[1705]) | ( l_46 [97] &  i[1705]);
assign l_45[50]    = ( l_46 [98] & !i[1705]) | ( l_46 [99] &  i[1705]);
assign l_45[51]    = ( l_46 [100] & !i[1705]) | ( l_46 [101] &  i[1705]);
assign l_45[52]    = ( l_46 [102] & !i[1705]) | ( l_46 [103] &  i[1705]);
assign l_45[53]    = ( l_46 [104] & !i[1705]) | ( l_46 [105] &  i[1705]);
assign l_45[54]    = ( l_46 [106] & !i[1705]) | ( l_46 [107] &  i[1705]);
assign l_45[55]    = ( l_46 [108] & !i[1705]) | ( l_46 [109] &  i[1705]);
assign l_45[56]    = ( l_46 [110] & !i[1705]) | ( l_46 [111] &  i[1705]);
assign l_45[57]    = ( l_46 [112] & !i[1705]) | ( l_46 [113] &  i[1705]);
assign l_45[58]    = ( l_46 [114] & !i[1705]) | ( l_46 [115] &  i[1705]);
assign l_45[59]    = ( l_46 [116] & !i[1705]) | ( l_46 [117] &  i[1705]);
assign l_45[60]    = ( l_46 [118] & !i[1705]) | ( l_46 [119] &  i[1705]);
assign l_45[61]    = ( l_46 [120] & !i[1705]) | ( l_46 [121] &  i[1705]);
assign l_45[62]    = ( l_46 [122] & !i[1705]) | ( l_46 [123] &  i[1705]);
assign l_45[63]    = ( l_46 [124] & !i[1705]) | ( l_46 [125] &  i[1705]);
assign l_45[64]    = ( l_46 [126] & !i[1705]) | ( l_46 [127] &  i[1705]);
assign l_45[65]    = ( l_46 [128] & !i[1705]) | ( l_46 [129] &  i[1705]);
assign l_45[66]    = ( l_46 [130] & !i[1705]) | ( l_46 [131] &  i[1705]);
assign l_45[67]    = ( l_46 [132] & !i[1705]) | ( l_46 [133] &  i[1705]);
assign l_45[68]    = ( l_46 [134] & !i[1705]) | ( l_46 [135] &  i[1705]);
assign l_45[69]    = ( l_46 [136] & !i[1705]) | ( l_46 [137] &  i[1705]);
assign l_45[70]    = ( l_46 [138] & !i[1705]) | ( l_46 [139] &  i[1705]);
assign l_45[71]    = ( l_46 [140] & !i[1705]) | ( l_46 [141] &  i[1705]);
assign l_45[72]    = ( l_46 [142] & !i[1705]) | ( l_46 [143] &  i[1705]);
assign l_45[73]    = ( l_46 [144] & !i[1705]) | ( l_46 [145] &  i[1705]);
assign l_45[74]    = ( l_46 [146] & !i[1705]) | ( l_46 [147] &  i[1705]);
assign l_45[75]    = ( l_46 [148] & !i[1705]) | ( l_46 [149] &  i[1705]);
assign l_45[76]    = ( l_46 [150] & !i[1705]) | ( l_46 [151] &  i[1705]);
assign l_45[77]    = ( l_46 [152] & !i[1705]) | ( l_46 [153] &  i[1705]);
assign l_45[78]    = ( l_46 [154] & !i[1705]) | ( l_46 [155] &  i[1705]);
assign l_45[79]    = ( l_46 [156] & !i[1705]) | ( l_46 [157] &  i[1705]);
assign l_45[80]    = ( l_46 [158] & !i[1705]) | ( l_46 [159] &  i[1705]);
assign l_45[81]    = ( l_46 [160] & !i[1705]) | ( l_46 [161] &  i[1705]);
assign l_45[82]    = ( l_46 [162] & !i[1705]) | ( l_46 [163] &  i[1705]);
assign l_45[83]    = ( l_46 [164] & !i[1705]) | ( l_46 [165] &  i[1705]);
assign l_45[84]    = ( l_46 [166] & !i[1705]) | ( l_46 [167] &  i[1705]);
assign l_45[85]    = ( l_46 [168] & !i[1705]) | ( l_46 [169] &  i[1705]);
assign l_45[86]    = ( l_46 [170] & !i[1705]) | ( l_46 [171] &  i[1705]);
assign l_45[87]    = ( l_46 [172] & !i[1705]) | ( l_46 [173] &  i[1705]);
assign l_45[88]    = ( l_46 [174] & !i[1705]) | ( l_46 [175] &  i[1705]);
assign l_45[89]    = ( l_46 [176] & !i[1705]) | ( l_46 [177] &  i[1705]);
assign l_45[90]    = ( l_46 [178] & !i[1705]) | ( l_46 [179] &  i[1705]);
assign l_45[91]    = ( l_46 [180] & !i[1705]) | ( l_46 [181] &  i[1705]);
assign l_45[92]    = ( l_46 [182] & !i[1705]) | ( l_46 [183] &  i[1705]);
assign l_45[93]    = ( l_46 [184] & !i[1705]) | ( l_46 [185] &  i[1705]);
assign l_45[94]    = ( l_46 [186] & !i[1705]) | ( l_46 [187] &  i[1705]);
assign l_45[95]    = ( l_46 [188] & !i[1705]) | ( l_46 [189] &  i[1705]);
assign l_45[96]    = ( l_46 [190] & !i[1705]) | ( l_46 [191] &  i[1705]);
assign l_45[97]    = ( l_46 [192] & !i[1705]) | ( l_46 [193] &  i[1705]);
assign l_45[98]    = ( l_46 [194] & !i[1705]) | ( l_46 [195] &  i[1705]);
assign l_45[99]    = ( l_46 [196] & !i[1705]) | ( l_46 [197] &  i[1705]);
assign l_45[100]    = ( l_46 [198] & !i[1705]) | ( l_46 [199] &  i[1705]);
assign l_45[101]    = ( l_46 [200] & !i[1705]) | ( l_46 [201] &  i[1705]);
assign l_45[102]    = ( l_46 [202] & !i[1705]) | ( l_46 [203] &  i[1705]);
assign l_45[103]    = ( l_46 [204] & !i[1705]) | ( l_46 [205] &  i[1705]);
assign l_45[104]    = ( l_46 [206] & !i[1705]) | ( l_46 [207] &  i[1705]);
assign l_45[105]    = ( l_46 [208] & !i[1705]) | ( l_46 [209] &  i[1705]);
assign l_45[106]    = ( l_46 [210] & !i[1705]) | ( l_46 [211] &  i[1705]);
assign l_45[107]    = ( l_46 [212] & !i[1705]) | ( l_46 [213] &  i[1705]);
assign l_45[108]    = ( l_46 [214] & !i[1705]) | ( l_46 [215] &  i[1705]);
assign l_45[109]    = ( l_46 [216] & !i[1705]) | ( l_46 [217] &  i[1705]);
assign l_45[110]    = ( l_46 [218] & !i[1705]) | ( l_46 [219] &  i[1705]);
assign l_45[111]    = ( l_46 [220] & !i[1705]) | ( l_46 [221] &  i[1705]);
assign l_45[112]    = ( l_46 [222] & !i[1705]) | ( l_46 [223] &  i[1705]);
assign l_45[113]    = ( l_46 [224] & !i[1705]) | ( l_46 [225] &  i[1705]);
assign l_45[114]    = ( l_46 [226] & !i[1705]) | ( l_46 [227] &  i[1705]);
assign l_45[115]    = ( l_46 [228] & !i[1705]) | ( l_46 [229] &  i[1705]);
assign l_45[116]    = ( l_46 [230] & !i[1705]) | ( l_46 [231] &  i[1705]);
assign l_45[117]    = ( l_46 [232] & !i[1705]) | ( l_46 [233] &  i[1705]);
assign l_45[118]    = ( l_46 [234] & !i[1705]) | ( l_46 [235] &  i[1705]);
assign l_45[119]    = ( l_46 [236] & !i[1705]) | ( l_46 [237] &  i[1705]);
assign l_45[120]    = ( l_46 [238] & !i[1705]) | ( l_46 [239] &  i[1705]);
assign l_45[121]    = ( l_46 [240] & !i[1705]) | ( l_46 [241] &  i[1705]);
assign l_45[122]    = ( l_46 [242] & !i[1705]) | ( l_46 [243] &  i[1705]);
assign l_45[123]    = ( l_46 [244] & !i[1705]) | ( l_46 [245] &  i[1705]);
assign l_45[124]    = ( l_46 [246] & !i[1705]) | ( l_46 [247] &  i[1705]);
assign l_45[125]    = ( l_46 [248] & !i[1705]) | ( l_46 [249] &  i[1705]);
assign l_45[126]    = ( l_46 [250] & !i[1705]) | ( l_46 [251] &  i[1705]);
assign l_45[127]    = ( l_46 [252] & !i[1705]) | ( l_46 [253] &  i[1705]);
assign l_45[128]    = ( l_46 [254] & !i[1705]) | ( l_46 [255] &  i[1705]);
assign l_45[129]    = ( l_46 [1] & !i[1705]) | ( l_46 [4] &  i[1705]);
assign l_45[130]    = ( l_46 [5] & !i[1705]) | ( l_46 [8] &  i[1705]);
assign l_45[131]    = ( l_46 [9] & !i[1705]) | ( l_46 [12] &  i[1705]);
assign l_45[132]    = ( l_46 [13] & !i[1705]) | ( l_46 [64] &  i[1705]);
assign l_45[133]    = ( l_46 [17] & !i[1705]) | ( l_46 [20] &  i[1705]);
assign l_45[134]    = ( l_46 [21] & !i[1705]) | ( l_46 [24] &  i[1705]);
assign l_45[135]    = ( l_46 [25] & !i[1705]) | ( l_46 [28] &  i[1705]);
assign l_45[136]    = ( l_46 [29] & !i[1705]) | ( l_46 [80] &  i[1705]);
assign l_45[137]    = ( l_46 [33] & !i[1705]) | ( l_46 [36] &  i[1705]);
assign l_45[138]    = ( l_46 [37] & !i[1705]) | ( l_46 [40] &  i[1705]);
assign l_45[139]    = ( l_46 [41] & !i[1705]) | ( l_46 [44] &  i[1705]);
assign l_45[140]    = ( l_46 [45] & !i[1705]) | ( l_46 [96] &  i[1705]);
assign l_45[141]    = ( l_46 [49] & !i[1705]) | ( l_46 [52] &  i[1705]);
assign l_45[142]    = ( l_46 [53] & !i[1705]) | ( l_46 [56] &  i[1705]);
assign l_45[143]    = ( l_46 [57] & !i[1705]) | ( l_46 [60] &  i[1705]);
assign l_45[144]    = ( l_46 [61] & !i[1705]) | ( l_46 [112] &  i[1705]);
assign l_45[145]    = ( l_46 [65] & !i[1705]) | ( l_46 [68] &  i[1705]);
assign l_45[146]    = ( l_46 [69] & !i[1705]) | ( l_46 [72] &  i[1705]);
assign l_45[147]    = ( l_46 [73] & !i[1705]) | ( l_46 [76] &  i[1705]);
assign l_45[148]    = ( l_46 [77] & !i[1705]) | ( l_46 [256] &  i[1705]);
assign l_45[149]    = ( l_46 [81] & !i[1705]) | ( l_46 [84] &  i[1705]);
assign l_45[150]    = ( l_46 [85] & !i[1705]) | ( l_46 [88] &  i[1705]);
assign l_45[151]    = ( l_46 [89] & !i[1705]) | ( l_46 [92] &  i[1705]);
assign l_45[152]    = ( l_46 [93] & !i[1705]) | ( l_46 [257] &  i[1705]);
assign l_45[153]    = ( l_46 [97] & !i[1705]) | ( l_46 [100] &  i[1705]);
assign l_45[154]    = ( l_46 [101] & !i[1705]) | ( l_46 [104] &  i[1705]);
assign l_45[155]    = ( l_46 [105] & !i[1705]) | ( l_46 [108] &  i[1705]);
assign l_45[156]    = ( l_46 [109] & !i[1705]) | ( l_46 [258] &  i[1705]);
assign l_45[157]    = ( l_46 [113] & !i[1705]) | ( l_46 [116] &  i[1705]);
assign l_45[158]    = ( l_46 [117] & !i[1705]) | ( l_46 [120] &  i[1705]);
assign l_45[159]    = ( l_46 [121] & !i[1705]) | ( l_46 [124] &  i[1705]);
assign l_45[160]    = ( l_46 [125] & !i[1705]) | ( l_46 [259] &  i[1705]);
assign l_45[161]    = ( l_46 [129] & !i[1705]) | ( l_46 [132] &  i[1705]);
assign l_45[162]    = ( l_46 [133] & !i[1705]) | ( l_46 [136] &  i[1705]);
assign l_45[163]    = ( l_46 [137] & !i[1705]) | ( l_46 [140] &  i[1705]);
assign l_45[164]    = ( l_46 [141] & !i[1705]) | ( l_46 [192] &  i[1705]);
assign l_45[165]    = ( l_46 [145] & !i[1705]) | ( l_46 [148] &  i[1705]);
assign l_45[166]    = ( l_46 [149] & !i[1705]) | ( l_46 [152] &  i[1705]);
assign l_45[167]    = ( l_46 [153] & !i[1705]) | ( l_46 [156] &  i[1705]);
assign l_45[168]    = ( l_46 [157] & !i[1705]) | ( l_46 [208] &  i[1705]);
assign l_45[169]    = ( l_46 [161] & !i[1705]) | ( l_46 [164] &  i[1705]);
assign l_45[170]    = ( l_46 [165] & !i[1705]) | ( l_46 [168] &  i[1705]);
assign l_45[171]    = ( l_46 [169] & !i[1705]) | ( l_46 [172] &  i[1705]);
assign l_45[172]    = ( l_46 [173] & !i[1705]) | ( l_46 [224] &  i[1705]);
assign l_45[173]    = ( l_46 [177] & !i[1705]) | ( l_46 [180] &  i[1705]);
assign l_45[174]    = ( l_46 [181] & !i[1705]) | ( l_46 [184] &  i[1705]);
assign l_45[175]    = ( l_46 [185] & !i[1705]) | ( l_46 [188] &  i[1705]);
assign l_45[176]    = ( l_46 [189] & !i[1705]) | ( l_46 [240] &  i[1705]);
assign l_45[177]    = ( l_46 [193] & !i[1705]) | ( l_46 [196] &  i[1705]);
assign l_45[178]    = ( l_46 [197] & !i[1705]) | ( l_46 [200] &  i[1705]);
assign l_45[179]    = ( l_46 [201] & !i[1705]) | ( l_46 [204] &  i[1705]);
assign l_45[180]    = ( l_46 [205] & !i[1705]) | ( l_46 [260] &  i[1705]);
assign l_45[181]    = ( l_46 [209] & !i[1705]) | ( l_46 [212] &  i[1705]);
assign l_45[182]    = ( l_46 [213] & !i[1705]) | ( l_46 [216] &  i[1705]);
assign l_45[183]    = ( l_46 [217] & !i[1705]) | ( l_46 [220] &  i[1705]);
assign l_45[184]    = ( l_46 [221] & !i[1705]) | ( l_46 [261] &  i[1705]);
assign l_45[185]    = ( l_46 [225] & !i[1705]) | ( l_46 [228] &  i[1705]);
assign l_45[186]    = ( l_46 [229] & !i[1705]) | ( l_46 [232] &  i[1705]);
assign l_45[187]    = ( l_46 [233] & !i[1705]) | ( l_46 [236] &  i[1705]);
assign l_45[188]    = ( l_46 [237] & !i[1705]) | ( l_46 [262] &  i[1705]);
assign l_45[189]    = ( l_46 [241] & !i[1705]) | ( l_46 [244] &  i[1705]);
assign l_45[190]    = ( l_46 [245] & !i[1705]) | ( l_46 [248] &  i[1705]);
assign l_45[191]    = ( l_46 [249] & !i[1705]) | ( l_46 [252] &  i[1705]);
assign l_45[192]    = ( l_46 [253] & !i[1705]) | ( l_46 [263] &  i[1705]);
assign l_45[193]    = ( l_46 [264] & !i[1705]) | ( l_46 [265] &  i[1705]);
assign l_45[194]    = ( l_46 [266] & !i[1705]) | ( l_46 [267] &  i[1705]);
assign l_45[195]    = ( l_46 [268] & !i[1705]) | ( l_46 [269] &  i[1705]);
assign l_45[196]    = ( l_46 [270] & !i[1705]) | ( l_46 [271] &  i[1705]);
assign l_45[197]    = ( l_46 [272] & !i[1705]) | ( l_46 [273] &  i[1705]);
assign l_45[198]    = ( l_46 [274] & !i[1705]) | ( l_46 [275] &  i[1705]);
assign l_45[199]    = ( l_46 [276] & !i[1705]) | ( l_46 [277] &  i[1705]);
assign l_45[200]    = ( l_46 [278] & !i[1705]) | ( l_46 [279] &  i[1705]);
assign l_45[201]    = ( l_46 [280] & !i[1705]) | ( l_46 [281] &  i[1705]);
assign l_45[202]    = ( l_46 [282] & !i[1705]) | ( l_46 [283] &  i[1705]);
assign l_45[203]    = ( l_46 [284] & !i[1705]) | ( l_46 [285] &  i[1705]);
assign l_45[204]    = ( l_46 [286] & !i[1705]) | ( l_46 [287] &  i[1705]);
assign l_45[205]    = ( l_46 [288] & !i[1705]) | ( l_46 [289] &  i[1705]);
assign l_45[206]    = ( l_46 [290] & !i[1705]) | ( l_46 [291] &  i[1705]);
assign l_45[207]    = ( l_46 [292] & !i[1705]) | ( l_46 [293] &  i[1705]);
assign l_45[208]    = ( l_46 [294] & !i[1705]) | ( l_46 [295] &  i[1705]);
assign l_45[209]    = ( l_46 [296] & !i[1705]) | ( l_46 [297] &  i[1705]);
assign l_45[210]    = ( l_46 [298] & !i[1705]) | ( l_46 [299] &  i[1705]);
assign l_45[211]    = ( l_46 [300] & !i[1705]) | ( l_46 [301] &  i[1705]);
assign l_45[212]    = ( l_46 [302] & !i[1705]) | ( l_46 [303] &  i[1705]);
assign l_45[213]    = ( l_46 [304] & !i[1705]) | ( l_46 [305] &  i[1705]);
assign l_45[214]    = ( l_46 [306] & !i[1705]) | ( l_46 [307] &  i[1705]);
assign l_45[215]    = ( l_46 [308] & !i[1705]) | ( l_46 [309] &  i[1705]);
assign l_45[216]    = ( l_46 [310] & !i[1705]) | ( l_46 [311] &  i[1705]);
assign l_45[217]    = ( l_46 [312] & !i[1705]) | ( l_46 [313] &  i[1705]);
assign l_45[218]    = ( l_46 [314] & !i[1705]) | ( l_46 [315] &  i[1705]);
assign l_45[219]    = ( l_46 [316] & !i[1705]) | ( l_46 [317] &  i[1705]);
assign l_45[220]    = ( l_46 [318] & !i[1705]) | ( l_46 [319] &  i[1705]);
assign l_45[221]    = ( l_46 [320] & !i[1705]) | ( l_46 [321] &  i[1705]);
assign l_45[222]    = ( l_46 [322] & !i[1705]) | ( l_46 [323] &  i[1705]);
assign l_45[223]    = ( l_46 [324] & !i[1705]) | ( l_46 [325] &  i[1705]);
assign l_45[224]    = ( l_46 [326] & !i[1705]) | ( l_46 [327] &  i[1705]);
assign l_45[225]    = ( l_46 [328]);
assign l_45[226]    = ( l_46 [329] & !i[1705]) | ( l_46 [330] &  i[1705]);
assign l_45[227]    = ( l_46 [331] & !i[1705]) | ( l_46 [332] &  i[1705]);
assign l_45[228]    = ( l_46 [333] & !i[1705]) | ( l_46 [334] &  i[1705]);
assign l_45[229]    = ( l_46 [335] & !i[1705]) | ( l_46 [336] &  i[1705]);
assign l_45[230]    = ( l_46 [337] & !i[1705]) | ( l_46 [338] &  i[1705]);
assign l_45[231]    = ( l_46 [339] & !i[1705]) | ( l_46 [340] &  i[1705]);
assign l_45[232]    = ( l_46 [341] & !i[1705]) | ( l_46 [342] &  i[1705]);
assign l_45[233]    = ( l_46 [343] & !i[1705]) | ( l_46 [344] &  i[1705]);
assign l_45[234]    = ( l_46 [345] & !i[1705]) | ( l_46 [346] &  i[1705]);
assign l_45[235]    = ( l_46 [347] & !i[1705]) | ( l_46 [348] &  i[1705]);
assign l_45[236]    = ( l_46 [349] & !i[1705]) | ( l_46 [350] &  i[1705]);
assign l_45[237]    = ( l_46 [351] & !i[1705]) | ( l_46 [352] &  i[1705]);
assign l_45[238]    = ( l_46 [353] & !i[1705]) | ( l_46 [354] &  i[1705]);
assign l_45[239]    = ( l_46 [355] & !i[1705]) | ( l_46 [356] &  i[1705]);
assign l_45[240]    = ( l_46 [357] & !i[1705]) | ( l_46 [358] &  i[1705]);
assign l_45[241]    = ( l_46 [359] & !i[1705]) | ( l_46 [360] &  i[1705]);
assign l_45[242]    = ( l_46 [361] & !i[1705]) | ( l_46 [362] &  i[1705]);
assign l_45[243]    = ( l_46 [363] & !i[1705]) | ( l_46 [364] &  i[1705]);
assign l_45[244]    = ( l_46 [365] & !i[1705]) | ( l_46 [366] &  i[1705]);
assign l_45[245]    = ( l_46 [367] & !i[1705]) | ( l_46 [368] &  i[1705]);
assign l_45[246]    = ( l_46 [369] & !i[1705]) | ( l_46 [370] &  i[1705]);
assign l_45[247]    = ( l_46 [371] & !i[1705]) | ( l_46 [372] &  i[1705]);
assign l_45[248]    = ( l_46 [373] & !i[1705]) | ( l_46 [374] &  i[1705]);
assign l_45[249]    = ( l_46 [375] & !i[1705]) | ( l_46 [376] &  i[1705]);
assign l_45[250]    = ( l_46 [377] & !i[1705]) | ( l_46 [378] &  i[1705]);
assign l_45[251]    = ( l_46 [379] & !i[1705]) | ( l_46 [380] &  i[1705]);
assign l_45[252]    = ( l_46 [381] & !i[1705]) | ( l_46 [382] &  i[1705]);
assign l_45[253]    = ( l_46 [383] & !i[1705]) | ( l_46 [384] &  i[1705]);
assign l_45[254]    = ( l_46 [385] & !i[1705]) | ( l_46 [386] &  i[1705]);
assign l_45[255]    = ( l_46 [387] & !i[1705]) | ( l_46 [388] &  i[1705]);
assign l_45[256]    = ( l_46 [389] & !i[1705]) | ( l_46 [390] &  i[1705]);
assign l_45[257]    = ( l_46 [391] & !i[1705]) | ( l_46 [392] &  i[1705]);
assign l_45[258]    = ( l_46 [393] & !i[1705]) | ( l_46 [394] &  i[1705]);
assign l_45[259]    = ( l_46 [395] & !i[1705]) | ( l_46 [396] &  i[1705]);
assign l_45[260]    = ( l_46 [397] & !i[1705]) | ( l_46 [398] &  i[1705]);
assign l_45[261]    = ( l_46 [399] & !i[1705]) | ( l_46 [400] &  i[1705]);
assign l_45[262]    = ( l_46 [401] & !i[1705]) | ( l_46 [402] &  i[1705]);
assign l_45[263]    = ( l_46 [403] & !i[1705]) | ( l_46 [404] &  i[1705]);
assign l_45[264]    = ( l_46 [405] & !i[1705]) | ( l_46 [406] &  i[1705]);
assign l_45[265]    = ( l_46 [407] & !i[1705]) | ( l_46 [408] &  i[1705]);
assign l_45[266]    = ( l_46 [409] & !i[1705]) | ( l_46 [410] &  i[1705]);
assign l_45[267]    = ( l_46 [411] & !i[1705]) | ( l_46 [412] &  i[1705]);
assign l_45[268]    = ( l_46 [413] & !i[1705]) | ( l_46 [414] &  i[1705]);
assign l_45[269]    = ( l_46 [415] & !i[1705]) | ( l_46 [416] &  i[1705]);
assign l_45[270]    = ( l_46 [417] & !i[1705]) | ( l_46 [418] &  i[1705]);
assign l_45[271]    = ( l_46 [419] & !i[1705]) | ( l_46 [420] &  i[1705]);
assign l_45[272]    = ( l_46 [421] & !i[1705]) | ( l_46 [422] &  i[1705]);
assign l_45[273]    = ( l_46 [423] & !i[1705]) | ( l_46 [424] &  i[1705]);
assign l_45[274]    = ( l_46 [425] & !i[1705]) | ( l_46 [426] &  i[1705]);
assign l_45[275]    = ( l_46 [427] & !i[1705]) | ( l_46 [428] &  i[1705]);
assign l_45[276]    = ( l_46 [429] & !i[1705]) | ( l_46 [430] &  i[1705]);
assign l_45[277]    = ( l_46 [431] & !i[1705]) | ( l_46 [432] &  i[1705]);
assign l_45[278]    = ( l_46 [433] & !i[1705]) | ( l_46 [434] &  i[1705]);
assign l_45[279]    = ( l_46 [435] & !i[1705]) | ( l_46 [436] &  i[1705]);
assign l_45[280]    = ( l_46 [437] & !i[1705]) | ( l_46 [438] &  i[1705]);
assign l_45[281]    = ( l_46 [439] & !i[1705]) | ( l_46 [440] &  i[1705]);
assign l_45[282]    = ( l_46 [441] & !i[1705]) | ( l_46 [442] &  i[1705]);
assign l_45[283]    = ( l_46 [443] & !i[1705]) | ( l_46 [444] &  i[1705]);
assign l_45[284]    = ( l_46 [445] & !i[1705]) | ( l_46 [446] &  i[1705]);
assign l_45[285]    = ( l_46 [447] & !i[1705]) | ( l_46 [448] &  i[1705]);
assign l_45[286]    = ( l_46 [449] & !i[1705]) | ( l_46 [450] &  i[1705]);
assign l_45[287]    = ( l_46 [451] & !i[1705]) | ( l_46 [452] &  i[1705]);
assign l_45[288]    = ( l_46 [453] & !i[1705]) | ( l_46 [454] &  i[1705]);
assign l_45[289]    = ( l_46 [455] & !i[1705]) | ( l_46 [456] &  i[1705]);
assign l_45[290]    = ( l_46 [457] & !i[1705]) | ( l_46 [458] &  i[1705]);
assign l_45[291]    = ( l_46 [459] & !i[1705]) | ( l_46 [460] &  i[1705]);
assign l_45[292]    = ( l_46 [461] & !i[1705]) | ( l_46 [462] &  i[1705]);
assign l_45[293]    = ( l_46 [463] & !i[1705]) | ( l_46 [464] &  i[1705]);
assign l_45[294]    = ( l_46 [465] & !i[1705]) | ( l_46 [466] &  i[1705]);
assign l_45[295]    = ( l_46 [467] & !i[1705]) | ( l_46 [468] &  i[1705]);
assign l_45[296]    = ( l_46 [469] & !i[1705]) | ( l_46 [470] &  i[1705]);
assign l_45[297]    = ( l_46 [471] & !i[1705]) | ( l_46 [472] &  i[1705]);
assign l_45[298]    = ( l_46 [473] & !i[1705]) | ( l_46 [474] &  i[1705]);
assign l_45[299]    = ( l_46 [475] & !i[1705]) | ( l_46 [476] &  i[1705]);
assign l_45[300]    = ( l_46 [477] & !i[1705]) | ( l_46 [478] &  i[1705]);
assign l_45[301]    = ( l_46 [479] & !i[1705]) | ( l_46 [480] &  i[1705]);
assign l_45[302]    = ( l_46 [481] & !i[1705]) | ( l_46 [482] &  i[1705]);
assign l_45[303]    = ( l_46 [483] & !i[1705]) | ( l_46 [484] &  i[1705]);
assign l_45[304]    = ( l_46 [485] & !i[1705]) | ( l_46 [486] &  i[1705]);
assign l_45[305]    = ( l_46 [487] & !i[1705]) | ( l_46 [488] &  i[1705]);
assign l_45[306]    = ( l_46 [489] & !i[1705]) | ( l_46 [490] &  i[1705]);
assign l_45[307]    = ( l_46 [491] & !i[1705]) | ( l_46 [492] &  i[1705]);
assign l_45[308]    = ( l_46 [493] & !i[1705]) | ( l_46 [494] &  i[1705]);
assign l_45[309]    = ( l_46 [495] & !i[1705]) | ( l_46 [496] &  i[1705]);
assign l_45[310]    = ( l_46 [497] & !i[1705]) | ( l_46 [498] &  i[1705]);
assign l_45[311]    = ( l_46 [499] & !i[1705]) | ( l_46 [500] &  i[1705]);
assign l_45[312]    = ( l_46 [501] & !i[1705]) | ( l_46 [502] &  i[1705]);
assign l_45[313]    = ( l_46 [503] & !i[1705]) | ( l_46 [504] &  i[1705]);
assign l_45[314]    = ( l_46 [505] & !i[1705]) | ( l_46 [506] &  i[1705]);
assign l_45[315]    = ( l_46 [507] & !i[1705]) | ( l_46 [508] &  i[1705]);
assign l_45[316]    = ( l_46 [509] & !i[1705]) | ( l_46 [510] &  i[1705]);
assign l_45[317]    = ( l_46 [511] & !i[1705]) | ( l_46 [512] &  i[1705]);
assign l_45[318]    = ( l_46 [513] & !i[1705]) | ( l_46 [514] &  i[1705]);
assign l_45[319]    = ( l_46 [515] & !i[1705]) | ( l_46 [516] &  i[1705]);
assign l_45[320]    = ( l_46 [517] & !i[1705]) | ( l_46 [518] &  i[1705]);
assign l_45[321]    = ( l_46 [519] & !i[1705]) | ( l_46 [520] &  i[1705]);
assign l_45[322]    = ( l_46 [265] & !i[1705]) | ( l_46 [268] &  i[1705]);
assign l_45[323]    = ( l_46 [269] & !i[1705]) | ( l_46 [272] &  i[1705]);
assign l_45[324]    = ( l_46 [273] & !i[1705]) | ( l_46 [276] &  i[1705]);
assign l_45[325]    = ( l_46 [277] & !i[1705]) | ( l_46 [329] &  i[1705]);
assign l_45[326]    = ( l_46 [281] & !i[1705]) | ( l_46 [284] &  i[1705]);
assign l_45[327]    = ( l_46 [285] & !i[1705]) | ( l_46 [288] &  i[1705]);
assign l_45[328]    = ( l_46 [289] & !i[1705]) | ( l_46 [292] &  i[1705]);
assign l_45[329]    = ( l_46 [293] & !i[1705]) | ( l_46 [345] &  i[1705]);
assign l_45[330]    = ( l_46 [297] & !i[1705]) | ( l_46 [300] &  i[1705]);
assign l_45[331]    = ( l_46 [301] & !i[1705]) | ( l_46 [304] &  i[1705]);
assign l_45[332]    = ( l_46 [305] & !i[1705]) | ( l_46 [308] &  i[1705]);
assign l_45[333]    = ( l_46 [309] & !i[1705]) | ( l_46 [361] &  i[1705]);
assign l_45[334]    = ( l_46 [313] & !i[1705]) | ( l_46 [316] &  i[1705]);
assign l_45[335]    = ( l_46 [317] & !i[1705]) | ( l_46 [320] &  i[1705]);
assign l_45[336]    = ( l_46 [321] & !i[1705]) | ( l_46 [324] &  i[1705]);
assign l_45[337]    = ( l_46 [325] & !i[1705]) | ( l_46 [377] &  i[1705]);
assign l_45[338]    = ( l_46 [330] & !i[1705]) | ( l_46 [333] &  i[1705]);
assign l_45[339]    = ( l_46 [334] & !i[1705]) | ( l_46 [337] &  i[1705]);
assign l_45[340]    = ( l_46 [338] & !i[1705]) | ( l_46 [341] &  i[1705]);
assign l_45[341]    = ( l_46 [342] & !i[1705]) | ( l_46 [521] &  i[1705]);
assign l_45[342]    = ( l_46 [346] & !i[1705]) | ( l_46 [349] &  i[1705]);
assign l_45[343]    = ( l_46 [350] & !i[1705]) | ( l_46 [353] &  i[1705]);
assign l_45[344]    = ( l_46 [354] & !i[1705]) | ( l_46 [357] &  i[1705]);
assign l_45[345]    = ( l_46 [358] & !i[1705]) | ( l_46 [522] &  i[1705]);
assign l_45[346]    = ( l_46 [362] & !i[1705]) | ( l_46 [365] &  i[1705]);
assign l_45[347]    = ( l_46 [366] & !i[1705]) | ( l_46 [369] &  i[1705]);
assign l_45[348]    = ( l_46 [370] & !i[1705]) | ( l_46 [373] &  i[1705]);
assign l_45[349]    = ( l_46 [374] & !i[1705]) | ( l_46 [523] &  i[1705]);
assign l_45[350]    = ( l_46 [378] & !i[1705]) | ( l_46 [381] &  i[1705]);
assign l_45[351]    = ( l_46 [382] & !i[1705]) | ( l_46 [385] &  i[1705]);
assign l_45[352]    = ( l_46 [386] & !i[1705]) | ( l_46 [389] &  i[1705]);
assign l_45[353]    = ( l_46 [390] & !i[1705]) | ( l_46 [524] &  i[1705]);
assign l_45[354]    = ( l_46 [394] & !i[1705]) | ( l_46 [397] &  i[1705]);
assign l_45[355]    = ( l_46 [398] & !i[1705]) | ( l_46 [401] &  i[1705]);
assign l_45[356]    = ( l_46 [402] & !i[1705]) | ( l_46 [405] &  i[1705]);
assign l_45[357]    = ( l_46 [406] & !i[1705]) | ( l_46 [457] &  i[1705]);
assign l_45[358]    = ( l_46 [410] & !i[1705]) | ( l_46 [413] &  i[1705]);
assign l_45[359]    = ( l_46 [414] & !i[1705]) | ( l_46 [417] &  i[1705]);
assign l_45[360]    = ( l_46 [418] & !i[1705]) | ( l_46 [421] &  i[1705]);
assign l_45[361]    = ( l_46 [422] & !i[1705]) | ( l_46 [473] &  i[1705]);
assign l_45[362]    = ( l_46 [426] & !i[1705]) | ( l_46 [429] &  i[1705]);
assign l_45[363]    = ( l_46 [430] & !i[1705]) | ( l_46 [433] &  i[1705]);
assign l_45[364]    = ( l_46 [434] & !i[1705]) | ( l_46 [437] &  i[1705]);
assign l_45[365]    = ( l_46 [438] & !i[1705]) | ( l_46 [489] &  i[1705]);
assign l_45[366]    = ( l_46 [442] & !i[1705]) | ( l_46 [445] &  i[1705]);
assign l_45[367]    = ( l_46 [446] & !i[1705]) | ( l_46 [449] &  i[1705]);
assign l_45[368]    = ( l_46 [450] & !i[1705]) | ( l_46 [453] &  i[1705]);
assign l_45[369]    = ( l_46 [454] & !i[1705]) | ( l_46 [505] &  i[1705]);
assign l_45[370]    = ( l_46 [458] & !i[1705]) | ( l_46 [461] &  i[1705]);
assign l_45[371]    = ( l_46 [462] & !i[1705]) | ( l_46 [465] &  i[1705]);
assign l_45[372]    = ( l_46 [466] & !i[1705]) | ( l_46 [469] &  i[1705]);
assign l_45[373]    = ( l_46 [470] & !i[1705]) | ( l_46 [525] &  i[1705]);
assign l_45[374]    = ( l_46 [474] & !i[1705]) | ( l_46 [477] &  i[1705]);
assign l_45[375]    = ( l_46 [478] & !i[1705]) | ( l_46 [481] &  i[1705]);
assign l_45[376]    = ( l_46 [482] & !i[1705]) | ( l_46 [485] &  i[1705]);
assign l_45[377]    = ( l_46 [486] & !i[1705]) | ( l_46 [526] &  i[1705]);
assign l_45[378]    = ( l_46 [490] & !i[1705]) | ( l_46 [493] &  i[1705]);
assign l_45[379]    = ( l_46 [494] & !i[1705]) | ( l_46 [497] &  i[1705]);
assign l_45[380]    = ( l_46 [498] & !i[1705]) | ( l_46 [501] &  i[1705]);
assign l_45[381]    = ( l_46 [502] & !i[1705]) | ( l_46 [527] &  i[1705]);
assign l_45[382]    = ( l_46 [506] & !i[1705]) | ( l_46 [509] &  i[1705]);
assign l_45[383]    = ( l_46 [510] & !i[1705]) | ( l_46 [513] &  i[1705]);
assign l_45[384]    = ( l_46 [514] & !i[1705]) | ( l_46 [517] &  i[1705]);
assign l_45[385]    = ( l_46 [518] & !i[1705]) | ( l_46 [528] &  i[1705]);
assign l_45[386]    = ( l_46 [529] &  i[1705]);
assign l_45[387]    = ( l_46 [530] & !i[1705]) | ( l_46 [531] &  i[1705]);
assign l_45[388]    = ( l_46 [532] & !i[1705]);
assign l_45[389]    = ( l_46 [532] & !i[1705]) | (      i[1705]);
assign l_45[390]    =  i[1705];
assign l_45[391]    = (!i[1705]) | ( l_46 [529] &  i[1705]);
assign l_45[392]    = ( l_46 [533] & !i[1705]) | ( l_46 [534] &  i[1705]);
assign l_45[393]    = ( l_46 [535] & !i[1705]) | ( l_46 [536] &  i[1705]);
assign l_46[0]    = ( l_47 [0] & !i[1821]) | ( l_47 [1] &  i[1821]);
assign l_46[1]    = ( l_47 [2] & !i[1821]) | ( l_47 [3] &  i[1821]);
assign l_46[2]    = ( l_47 [4] & !i[1821]) | ( l_47 [5] &  i[1821]);
assign l_46[3]    = ( l_47 [6] & !i[1821]) | ( l_47 [7] &  i[1821]);
assign l_46[4]    = ( l_47 [8] & !i[1821]) | ( l_47 [9] &  i[1821]);
assign l_46[5]    = ( l_47 [10] & !i[1821]) | ( l_47 [11] &  i[1821]);
assign l_46[6]    = ( l_47 [12] & !i[1821]) | ( l_47 [13] &  i[1821]);
assign l_46[7]    = ( l_47 [14] & !i[1821]) | ( l_47 [15] &  i[1821]);
assign l_46[8]    = ( l_47 [16] & !i[1821]) | ( l_47 [17] &  i[1821]);
assign l_46[9]    = ( l_47 [18] & !i[1821]) | ( l_47 [19] &  i[1821]);
assign l_46[10]    = ( l_47 [20] & !i[1821]) | ( l_47 [21] &  i[1821]);
assign l_46[11]    = ( l_47 [22] & !i[1821]) | ( l_47 [23] &  i[1821]);
assign l_46[12]    = ( l_47 [24] & !i[1821]) | ( l_47 [25] &  i[1821]);
assign l_46[13]    = ( l_47 [26] & !i[1821]) | ( l_47 [27] &  i[1821]);
assign l_46[14]    = ( l_47 [28] & !i[1821]) | ( l_47 [29] &  i[1821]);
assign l_46[15]    = ( l_47 [30] & !i[1821]) | ( l_47 [31] &  i[1821]);
assign l_46[16]    = ( l_47 [32] & !i[1821]) | ( l_47 [33] &  i[1821]);
assign l_46[17]    = ( l_47 [34] & !i[1821]) | ( l_47 [35] &  i[1821]);
assign l_46[18]    = ( l_47 [36] & !i[1821]) | ( l_47 [37] &  i[1821]);
assign l_46[19]    = ( l_47 [38] & !i[1821]) | ( l_47 [39] &  i[1821]);
assign l_46[20]    = ( l_47 [40] & !i[1821]) | ( l_47 [41] &  i[1821]);
assign l_46[21]    = ( l_47 [42] & !i[1821]) | ( l_47 [43] &  i[1821]);
assign l_46[22]    = ( l_47 [44] & !i[1821]) | ( l_47 [45] &  i[1821]);
assign l_46[23]    = ( l_47 [46] & !i[1821]) | ( l_47 [47] &  i[1821]);
assign l_46[24]    = ( l_47 [48] & !i[1821]) | ( l_47 [49] &  i[1821]);
assign l_46[25]    = ( l_47 [50] & !i[1821]) | ( l_47 [51] &  i[1821]);
assign l_46[26]    = ( l_47 [52] & !i[1821]) | ( l_47 [53] &  i[1821]);
assign l_46[27]    = ( l_47 [54] & !i[1821]) | ( l_47 [55] &  i[1821]);
assign l_46[28]    = ( l_47 [56] & !i[1821]) | ( l_47 [57] &  i[1821]);
assign l_46[29]    = ( l_47 [58] & !i[1821]) | ( l_47 [59] &  i[1821]);
assign l_46[30]    = ( l_47 [60] & !i[1821]) | ( l_47 [61] &  i[1821]);
assign l_46[31]    = ( l_47 [62] & !i[1821]) | ( l_47 [63] &  i[1821]);
assign l_46[32]    = ( l_47 [64] & !i[1821]) | ( l_47 [65] &  i[1821]);
assign l_46[33]    = ( l_47 [66] & !i[1821]) | ( l_47 [67] &  i[1821]);
assign l_46[34]    = ( l_47 [68] & !i[1821]) | ( l_47 [69] &  i[1821]);
assign l_46[35]    = ( l_47 [70] & !i[1821]) | ( l_47 [71] &  i[1821]);
assign l_46[36]    = ( l_47 [72] & !i[1821]) | ( l_47 [73] &  i[1821]);
assign l_46[37]    = ( l_47 [74] & !i[1821]) | ( l_47 [75] &  i[1821]);
assign l_46[38]    = ( l_47 [76] & !i[1821]) | ( l_47 [77] &  i[1821]);
assign l_46[39]    = ( l_47 [78] & !i[1821]) | ( l_47 [79] &  i[1821]);
assign l_46[40]    = ( l_47 [80] & !i[1821]) | ( l_47 [81] &  i[1821]);
assign l_46[41]    = ( l_47 [82] & !i[1821]) | ( l_47 [83] &  i[1821]);
assign l_46[42]    = ( l_47 [84] & !i[1821]) | ( l_47 [85] &  i[1821]);
assign l_46[43]    = ( l_47 [86] & !i[1821]) | ( l_47 [87] &  i[1821]);
assign l_46[44]    = ( l_47 [88] & !i[1821]) | ( l_47 [89] &  i[1821]);
assign l_46[45]    = ( l_47 [90] & !i[1821]) | ( l_47 [91] &  i[1821]);
assign l_46[46]    = ( l_47 [92] & !i[1821]) | ( l_47 [93] &  i[1821]);
assign l_46[47]    = ( l_47 [94] & !i[1821]) | ( l_47 [95] &  i[1821]);
assign l_46[48]    = ( l_47 [96] & !i[1821]) | ( l_47 [97] &  i[1821]);
assign l_46[49]    = ( l_47 [98] & !i[1821]) | ( l_47 [99] &  i[1821]);
assign l_46[50]    = ( l_47 [100] & !i[1821]) | ( l_47 [101] &  i[1821]);
assign l_46[51]    = ( l_47 [102] & !i[1821]) | ( l_47 [103] &  i[1821]);
assign l_46[52]    = ( l_47 [104] & !i[1821]) | ( l_47 [105] &  i[1821]);
assign l_46[53]    = ( l_47 [106] & !i[1821]) | ( l_47 [107] &  i[1821]);
assign l_46[54]    = ( l_47 [108] & !i[1821]) | ( l_47 [109] &  i[1821]);
assign l_46[55]    = ( l_47 [110] & !i[1821]) | ( l_47 [111] &  i[1821]);
assign l_46[56]    = ( l_47 [112] & !i[1821]) | ( l_47 [113] &  i[1821]);
assign l_46[57]    = ( l_47 [114] & !i[1821]) | ( l_47 [115] &  i[1821]);
assign l_46[58]    = ( l_47 [116] & !i[1821]) | ( l_47 [117] &  i[1821]);
assign l_46[59]    = ( l_47 [118] & !i[1821]) | ( l_47 [119] &  i[1821]);
assign l_46[60]    = ( l_47 [120] & !i[1821]) | ( l_47 [121] &  i[1821]);
assign l_46[61]    = ( l_47 [122] & !i[1821]) | ( l_47 [123] &  i[1821]);
assign l_46[62]    = ( l_47 [124] & !i[1821]) | ( l_47 [125] &  i[1821]);
assign l_46[63]    = ( l_47 [126] & !i[1821]) | ( l_47 [127] &  i[1821]);
assign l_46[64]    = ( l_47 [128] & !i[1821]) | ( l_47 [129] &  i[1821]);
assign l_46[65]    = ( l_47 [130] & !i[1821]) | ( l_47 [131] &  i[1821]);
assign l_46[66]    = ( l_47 [132] & !i[1821]) | ( l_47 [133] &  i[1821]);
assign l_46[67]    = ( l_47 [134] & !i[1821]) | ( l_47 [135] &  i[1821]);
assign l_46[68]    = ( l_47 [136] & !i[1821]) | ( l_47 [137] &  i[1821]);
assign l_46[69]    = ( l_47 [138] & !i[1821]) | ( l_47 [139] &  i[1821]);
assign l_46[70]    = ( l_47 [140] & !i[1821]) | ( l_47 [141] &  i[1821]);
assign l_46[71]    = ( l_47 [142] & !i[1821]) | ( l_47 [143] &  i[1821]);
assign l_46[72]    = ( l_47 [144] & !i[1821]) | ( l_47 [145] &  i[1821]);
assign l_46[73]    = ( l_47 [146] & !i[1821]) | ( l_47 [147] &  i[1821]);
assign l_46[74]    = ( l_47 [148] & !i[1821]) | ( l_47 [149] &  i[1821]);
assign l_46[75]    = ( l_47 [150] & !i[1821]) | ( l_47 [151] &  i[1821]);
assign l_46[76]    = ( l_47 [152] & !i[1821]) | ( l_47 [153] &  i[1821]);
assign l_46[77]    = ( l_47 [154] & !i[1821]) | ( l_47 [155] &  i[1821]);
assign l_46[78]    = ( l_47 [156] & !i[1821]) | ( l_47 [157] &  i[1821]);
assign l_46[79]    = ( l_47 [158] & !i[1821]) | ( l_47 [159] &  i[1821]);
assign l_46[80]    = ( l_47 [160] & !i[1821]) | ( l_47 [161] &  i[1821]);
assign l_46[81]    = ( l_47 [162] & !i[1821]) | ( l_47 [163] &  i[1821]);
assign l_46[82]    = ( l_47 [164] & !i[1821]) | ( l_47 [165] &  i[1821]);
assign l_46[83]    = ( l_47 [166] & !i[1821]) | ( l_47 [167] &  i[1821]);
assign l_46[84]    = ( l_47 [168] & !i[1821]) | ( l_47 [169] &  i[1821]);
assign l_46[85]    = ( l_47 [170] & !i[1821]) | ( l_47 [171] &  i[1821]);
assign l_46[86]    = ( l_47 [172] & !i[1821]) | ( l_47 [173] &  i[1821]);
assign l_46[87]    = ( l_47 [174] & !i[1821]) | ( l_47 [175] &  i[1821]);
assign l_46[88]    = ( l_47 [176] & !i[1821]) | ( l_47 [177] &  i[1821]);
assign l_46[89]    = ( l_47 [178] & !i[1821]) | ( l_47 [179] &  i[1821]);
assign l_46[90]    = ( l_47 [180] & !i[1821]) | ( l_47 [181] &  i[1821]);
assign l_46[91]    = ( l_47 [182] & !i[1821]) | ( l_47 [183] &  i[1821]);
assign l_46[92]    = ( l_47 [184] & !i[1821]) | ( l_47 [185] &  i[1821]);
assign l_46[93]    = ( l_47 [186] & !i[1821]) | ( l_47 [187] &  i[1821]);
assign l_46[94]    = ( l_47 [188] & !i[1821]) | ( l_47 [189] &  i[1821]);
assign l_46[95]    = ( l_47 [190] & !i[1821]) | ( l_47 [191] &  i[1821]);
assign l_46[96]    = ( l_47 [192] & !i[1821]) | ( l_47 [193] &  i[1821]);
assign l_46[97]    = ( l_47 [194] & !i[1821]) | ( l_47 [195] &  i[1821]);
assign l_46[98]    = ( l_47 [196] & !i[1821]) | ( l_47 [197] &  i[1821]);
assign l_46[99]    = ( l_47 [198] & !i[1821]) | ( l_47 [199] &  i[1821]);
assign l_46[100]    = ( l_47 [200] & !i[1821]) | ( l_47 [201] &  i[1821]);
assign l_46[101]    = ( l_47 [202] & !i[1821]) | ( l_47 [203] &  i[1821]);
assign l_46[102]    = ( l_47 [204] & !i[1821]) | ( l_47 [205] &  i[1821]);
assign l_46[103]    = ( l_47 [206] & !i[1821]) | ( l_47 [207] &  i[1821]);
assign l_46[104]    = ( l_47 [208] & !i[1821]) | ( l_47 [209] &  i[1821]);
assign l_46[105]    = ( l_47 [210] & !i[1821]) | ( l_47 [211] &  i[1821]);
assign l_46[106]    = ( l_47 [212] & !i[1821]) | ( l_47 [213] &  i[1821]);
assign l_46[107]    = ( l_47 [214] & !i[1821]) | ( l_47 [215] &  i[1821]);
assign l_46[108]    = ( l_47 [216] & !i[1821]) | ( l_47 [217] &  i[1821]);
assign l_46[109]    = ( l_47 [218] & !i[1821]) | ( l_47 [219] &  i[1821]);
assign l_46[110]    = ( l_47 [220] & !i[1821]) | ( l_47 [221] &  i[1821]);
assign l_46[111]    = ( l_47 [222] & !i[1821]) | ( l_47 [223] &  i[1821]);
assign l_46[112]    = ( l_47 [224] & !i[1821]) | ( l_47 [225] &  i[1821]);
assign l_46[113]    = ( l_47 [226] & !i[1821]) | ( l_47 [227] &  i[1821]);
assign l_46[114]    = ( l_47 [228] & !i[1821]) | ( l_47 [229] &  i[1821]);
assign l_46[115]    = ( l_47 [230] & !i[1821]) | ( l_47 [231] &  i[1821]);
assign l_46[116]    = ( l_47 [232] & !i[1821]) | ( l_47 [233] &  i[1821]);
assign l_46[117]    = ( l_47 [234] & !i[1821]) | ( l_47 [235] &  i[1821]);
assign l_46[118]    = ( l_47 [236] & !i[1821]) | ( l_47 [237] &  i[1821]);
assign l_46[119]    = ( l_47 [238] & !i[1821]) | ( l_47 [239] &  i[1821]);
assign l_46[120]    = ( l_47 [240] & !i[1821]) | ( l_47 [241] &  i[1821]);
assign l_46[121]    = ( l_47 [242] & !i[1821]) | ( l_47 [243] &  i[1821]);
assign l_46[122]    = ( l_47 [244] & !i[1821]) | ( l_47 [245] &  i[1821]);
assign l_46[123]    = ( l_47 [246] & !i[1821]) | ( l_47 [247] &  i[1821]);
assign l_46[124]    = ( l_47 [248] & !i[1821]) | ( l_47 [249] &  i[1821]);
assign l_46[125]    = ( l_47 [250] & !i[1821]) | ( l_47 [251] &  i[1821]);
assign l_46[126]    = ( l_47 [252] & !i[1821]) | ( l_47 [253] &  i[1821]);
assign l_46[127]    = ( l_47 [254] & !i[1821]) | ( l_47 [255] &  i[1821]);
assign l_46[128]    = ( l_47 [256] & !i[1821]) | ( l_47 [257] &  i[1821]);
assign l_46[129]    = ( l_47 [258] & !i[1821]) | ( l_47 [259] &  i[1821]);
assign l_46[130]    = ( l_47 [260] & !i[1821]) | ( l_47 [261] &  i[1821]);
assign l_46[131]    = ( l_47 [262] & !i[1821]) | ( l_47 [263] &  i[1821]);
assign l_46[132]    = ( l_47 [264] & !i[1821]) | ( l_47 [265] &  i[1821]);
assign l_46[133]    = ( l_47 [266] & !i[1821]) | ( l_47 [267] &  i[1821]);
assign l_46[134]    = ( l_47 [268] & !i[1821]) | ( l_47 [269] &  i[1821]);
assign l_46[135]    = ( l_47 [270] & !i[1821]) | ( l_47 [271] &  i[1821]);
assign l_46[136]    = ( l_47 [272] & !i[1821]) | ( l_47 [273] &  i[1821]);
assign l_46[137]    = ( l_47 [274] & !i[1821]) | ( l_47 [275] &  i[1821]);
assign l_46[138]    = ( l_47 [276] & !i[1821]) | ( l_47 [277] &  i[1821]);
assign l_46[139]    = ( l_47 [278] & !i[1821]) | ( l_47 [279] &  i[1821]);
assign l_46[140]    = ( l_47 [280] & !i[1821]) | ( l_47 [281] &  i[1821]);
assign l_46[141]    = ( l_47 [282] & !i[1821]) | ( l_47 [283] &  i[1821]);
assign l_46[142]    = ( l_47 [284] & !i[1821]) | ( l_47 [285] &  i[1821]);
assign l_46[143]    = ( l_47 [286] & !i[1821]) | ( l_47 [287] &  i[1821]);
assign l_46[144]    = ( l_47 [288] & !i[1821]) | ( l_47 [289] &  i[1821]);
assign l_46[145]    = ( l_47 [290] & !i[1821]) | ( l_47 [291] &  i[1821]);
assign l_46[146]    = ( l_47 [292] & !i[1821]) | ( l_47 [293] &  i[1821]);
assign l_46[147]    = ( l_47 [294] & !i[1821]) | ( l_47 [295] &  i[1821]);
assign l_46[148]    = ( l_47 [296] & !i[1821]) | ( l_47 [297] &  i[1821]);
assign l_46[149]    = ( l_47 [298] & !i[1821]) | ( l_47 [299] &  i[1821]);
assign l_46[150]    = ( l_47 [300] & !i[1821]) | ( l_47 [301] &  i[1821]);
assign l_46[151]    = ( l_47 [302] & !i[1821]) | ( l_47 [303] &  i[1821]);
assign l_46[152]    = ( l_47 [304] & !i[1821]) | ( l_47 [305] &  i[1821]);
assign l_46[153]    = ( l_47 [306] & !i[1821]) | ( l_47 [307] &  i[1821]);
assign l_46[154]    = ( l_47 [308] & !i[1821]) | ( l_47 [309] &  i[1821]);
assign l_46[155]    = ( l_47 [310] & !i[1821]) | ( l_47 [311] &  i[1821]);
assign l_46[156]    = ( l_47 [312] & !i[1821]) | ( l_47 [313] &  i[1821]);
assign l_46[157]    = ( l_47 [314] & !i[1821]) | ( l_47 [315] &  i[1821]);
assign l_46[158]    = ( l_47 [316] & !i[1821]) | ( l_47 [317] &  i[1821]);
assign l_46[159]    = ( l_47 [318] & !i[1821]) | ( l_47 [319] &  i[1821]);
assign l_46[160]    = ( l_47 [320] & !i[1821]) | ( l_47 [321] &  i[1821]);
assign l_46[161]    = ( l_47 [322] & !i[1821]) | ( l_47 [323] &  i[1821]);
assign l_46[162]    = ( l_47 [324] & !i[1821]) | ( l_47 [325] &  i[1821]);
assign l_46[163]    = ( l_47 [326] & !i[1821]) | ( l_47 [327] &  i[1821]);
assign l_46[164]    = ( l_47 [328] & !i[1821]) | ( l_47 [329] &  i[1821]);
assign l_46[165]    = ( l_47 [330] & !i[1821]) | ( l_47 [331] &  i[1821]);
assign l_46[166]    = ( l_47 [332] & !i[1821]) | ( l_47 [333] &  i[1821]);
assign l_46[167]    = ( l_47 [334] & !i[1821]) | ( l_47 [335] &  i[1821]);
assign l_46[168]    = ( l_47 [336] & !i[1821]) | ( l_47 [337] &  i[1821]);
assign l_46[169]    = ( l_47 [338] & !i[1821]) | ( l_47 [339] &  i[1821]);
assign l_46[170]    = ( l_47 [340] & !i[1821]) | ( l_47 [341] &  i[1821]);
assign l_46[171]    = ( l_47 [342] & !i[1821]) | ( l_47 [343] &  i[1821]);
assign l_46[172]    = ( l_47 [344] & !i[1821]) | ( l_47 [345] &  i[1821]);
assign l_46[173]    = ( l_47 [346] & !i[1821]) | ( l_47 [347] &  i[1821]);
assign l_46[174]    = ( l_47 [348] & !i[1821]) | ( l_47 [349] &  i[1821]);
assign l_46[175]    = ( l_47 [350] & !i[1821]) | ( l_47 [351] &  i[1821]);
assign l_46[176]    = ( l_47 [352] & !i[1821]) | ( l_47 [353] &  i[1821]);
assign l_46[177]    = ( l_47 [354] & !i[1821]) | ( l_47 [355] &  i[1821]);
assign l_46[178]    = ( l_47 [356] & !i[1821]) | ( l_47 [357] &  i[1821]);
assign l_46[179]    = ( l_47 [358] & !i[1821]) | ( l_47 [359] &  i[1821]);
assign l_46[180]    = ( l_47 [360] & !i[1821]) | ( l_47 [361] &  i[1821]);
assign l_46[181]    = ( l_47 [362] & !i[1821]) | ( l_47 [363] &  i[1821]);
assign l_46[182]    = ( l_47 [364] & !i[1821]) | ( l_47 [365] &  i[1821]);
assign l_46[183]    = ( l_47 [366] & !i[1821]) | ( l_47 [367] &  i[1821]);
assign l_46[184]    = ( l_47 [368] & !i[1821]) | ( l_47 [369] &  i[1821]);
assign l_46[185]    = ( l_47 [370] & !i[1821]) | ( l_47 [371] &  i[1821]);
assign l_46[186]    = ( l_47 [372] & !i[1821]) | ( l_47 [373] &  i[1821]);
assign l_46[187]    = ( l_47 [374] & !i[1821]) | ( l_47 [375] &  i[1821]);
assign l_46[188]    = ( l_47 [376] & !i[1821]) | ( l_47 [377] &  i[1821]);
assign l_46[189]    = ( l_47 [378] & !i[1821]) | ( l_47 [379] &  i[1821]);
assign l_46[190]    = ( l_47 [380] & !i[1821]) | ( l_47 [381] &  i[1821]);
assign l_46[191]    = ( l_47 [382] & !i[1821]) | ( l_47 [383] &  i[1821]);
assign l_46[192]    = ( l_47 [384] & !i[1821]) | ( l_47 [385] &  i[1821]);
assign l_46[193]    = ( l_47 [386] & !i[1821]) | ( l_47 [387] &  i[1821]);
assign l_46[194]    = ( l_47 [388] & !i[1821]) | ( l_47 [389] &  i[1821]);
assign l_46[195]    = ( l_47 [390] & !i[1821]) | ( l_47 [391] &  i[1821]);
assign l_46[196]    = ( l_47 [392] & !i[1821]) | ( l_47 [393] &  i[1821]);
assign l_46[197]    = ( l_47 [394] & !i[1821]) | ( l_47 [395] &  i[1821]);
assign l_46[198]    = ( l_47 [396] & !i[1821]) | ( l_47 [397] &  i[1821]);
assign l_46[199]    = ( l_47 [398] & !i[1821]) | ( l_47 [399] &  i[1821]);
assign l_46[200]    = ( l_47 [400] & !i[1821]) | ( l_47 [401] &  i[1821]);
assign l_46[201]    = ( l_47 [402] & !i[1821]) | ( l_47 [403] &  i[1821]);
assign l_46[202]    = ( l_47 [404] & !i[1821]) | ( l_47 [405] &  i[1821]);
assign l_46[203]    = ( l_47 [406] & !i[1821]) | ( l_47 [407] &  i[1821]);
assign l_46[204]    = ( l_47 [408] & !i[1821]) | ( l_47 [409] &  i[1821]);
assign l_46[205]    = ( l_47 [410] & !i[1821]) | ( l_47 [411] &  i[1821]);
assign l_46[206]    = ( l_47 [412] & !i[1821]) | ( l_47 [413] &  i[1821]);
assign l_46[207]    = ( l_47 [414] & !i[1821]) | ( l_47 [415] &  i[1821]);
assign l_46[208]    = ( l_47 [416] & !i[1821]) | ( l_47 [417] &  i[1821]);
assign l_46[209]    = ( l_47 [418] & !i[1821]) | ( l_47 [419] &  i[1821]);
assign l_46[210]    = ( l_47 [420] & !i[1821]) | ( l_47 [421] &  i[1821]);
assign l_46[211]    = ( l_47 [422] & !i[1821]) | ( l_47 [423] &  i[1821]);
assign l_46[212]    = ( l_47 [424] & !i[1821]) | ( l_47 [425] &  i[1821]);
assign l_46[213]    = ( l_47 [426] & !i[1821]) | ( l_47 [427] &  i[1821]);
assign l_46[214]    = ( l_47 [428] & !i[1821]) | ( l_47 [429] &  i[1821]);
assign l_46[215]    = ( l_47 [430] & !i[1821]) | ( l_47 [431] &  i[1821]);
assign l_46[216]    = ( l_47 [432] & !i[1821]) | ( l_47 [433] &  i[1821]);
assign l_46[217]    = ( l_47 [434] & !i[1821]) | ( l_47 [435] &  i[1821]);
assign l_46[218]    = ( l_47 [436] & !i[1821]) | ( l_47 [437] &  i[1821]);
assign l_46[219]    = ( l_47 [438] & !i[1821]) | ( l_47 [439] &  i[1821]);
assign l_46[220]    = ( l_47 [440] & !i[1821]) | ( l_47 [441] &  i[1821]);
assign l_46[221]    = ( l_47 [442] & !i[1821]) | ( l_47 [443] &  i[1821]);
assign l_46[222]    = ( l_47 [444] & !i[1821]) | ( l_47 [445] &  i[1821]);
assign l_46[223]    = ( l_47 [446] & !i[1821]) | ( l_47 [447] &  i[1821]);
assign l_46[224]    = ( l_47 [448] & !i[1821]) | ( l_47 [449] &  i[1821]);
assign l_46[225]    = ( l_47 [450] & !i[1821]) | ( l_47 [451] &  i[1821]);
assign l_46[226]    = ( l_47 [452] & !i[1821]) | ( l_47 [453] &  i[1821]);
assign l_46[227]    = ( l_47 [454] & !i[1821]) | ( l_47 [455] &  i[1821]);
assign l_46[228]    = ( l_47 [456] & !i[1821]) | ( l_47 [457] &  i[1821]);
assign l_46[229]    = ( l_47 [458] & !i[1821]) | ( l_47 [459] &  i[1821]);
assign l_46[230]    = ( l_47 [460] & !i[1821]) | ( l_47 [461] &  i[1821]);
assign l_46[231]    = ( l_47 [462] & !i[1821]) | ( l_47 [463] &  i[1821]);
assign l_46[232]    = ( l_47 [464] & !i[1821]) | ( l_47 [465] &  i[1821]);
assign l_46[233]    = ( l_47 [466] & !i[1821]) | ( l_47 [467] &  i[1821]);
assign l_46[234]    = ( l_47 [468] & !i[1821]) | ( l_47 [469] &  i[1821]);
assign l_46[235]    = ( l_47 [470] & !i[1821]) | ( l_47 [471] &  i[1821]);
assign l_46[236]    = ( l_47 [472] & !i[1821]) | ( l_47 [473] &  i[1821]);
assign l_46[237]    = ( l_47 [474] & !i[1821]) | ( l_47 [475] &  i[1821]);
assign l_46[238]    = ( l_47 [476] & !i[1821]) | ( l_47 [477] &  i[1821]);
assign l_46[239]    = ( l_47 [478] & !i[1821]) | ( l_47 [479] &  i[1821]);
assign l_46[240]    = ( l_47 [480] & !i[1821]) | ( l_47 [481] &  i[1821]);
assign l_46[241]    = ( l_47 [482] & !i[1821]) | ( l_47 [483] &  i[1821]);
assign l_46[242]    = ( l_47 [484] & !i[1821]) | ( l_47 [485] &  i[1821]);
assign l_46[243]    = ( l_47 [486] & !i[1821]) | ( l_47 [487] &  i[1821]);
assign l_46[244]    = ( l_47 [488] & !i[1821]) | ( l_47 [489] &  i[1821]);
assign l_46[245]    = ( l_47 [490] & !i[1821]) | ( l_47 [491] &  i[1821]);
assign l_46[246]    = ( l_47 [492] & !i[1821]) | ( l_47 [493] &  i[1821]);
assign l_46[247]    = ( l_47 [494] & !i[1821]) | ( l_47 [495] &  i[1821]);
assign l_46[248]    = ( l_47 [496] & !i[1821]) | ( l_47 [497] &  i[1821]);
assign l_46[249]    = ( l_47 [498] & !i[1821]) | ( l_47 [499] &  i[1821]);
assign l_46[250]    = ( l_47 [500] & !i[1821]) | ( l_47 [501] &  i[1821]);
assign l_46[251]    = ( l_47 [502] & !i[1821]) | ( l_47 [503] &  i[1821]);
assign l_46[252]    = ( l_47 [504] & !i[1821]) | ( l_47 [505] &  i[1821]);
assign l_46[253]    = ( l_47 [506] & !i[1821]) | ( l_47 [507] &  i[1821]);
assign l_46[254]    = ( l_47 [508] & !i[1821]) | ( l_47 [509] &  i[1821]);
assign l_46[255]    = ( l_47 [510] & !i[1821]) | ( l_47 [511] &  i[1821]);
assign l_46[256]    = ( l_47 [512] & !i[1821]) | ( l_47 [513] &  i[1821]);
assign l_46[257]    = ( l_47 [514] & !i[1821]) | ( l_47 [515] &  i[1821]);
assign l_46[258]    = ( l_47 [516] & !i[1821]) | ( l_47 [517] &  i[1821]);
assign l_46[259]    = ( l_47 [518] & !i[1821]) | ( l_47 [519] &  i[1821]);
assign l_46[260]    = ( l_47 [520] & !i[1821]) | ( l_47 [521] &  i[1821]);
assign l_46[261]    = ( l_47 [522] & !i[1821]) | ( l_47 [523] &  i[1821]);
assign l_46[262]    = ( l_47 [524] & !i[1821]) | ( l_47 [525] &  i[1821]);
assign l_46[263]    = ( l_47 [526] & !i[1821]) | ( l_47 [527] &  i[1821]);
assign l_46[264]    = ( l_47 [528] & !i[1821]) | ( l_47 [529] &  i[1821]);
assign l_46[265]    = ( l_47 [530] & !i[1821]) | ( l_47 [531] &  i[1821]);
assign l_46[266]    = ( l_47 [532] & !i[1821]) | ( l_47 [533] &  i[1821]);
assign l_46[267]    = ( l_47 [534] & !i[1821]) | ( l_47 [535] &  i[1821]);
assign l_46[268]    = ( l_47 [536] & !i[1821]) | ( l_47 [537] &  i[1821]);
assign l_46[269]    = ( l_47 [538] & !i[1821]) | ( l_47 [539] &  i[1821]);
assign l_46[270]    = ( l_47 [540] & !i[1821]) | ( l_47 [541] &  i[1821]);
assign l_46[271]    = ( l_47 [542] & !i[1821]) | ( l_47 [543] &  i[1821]);
assign l_46[272]    = ( l_47 [544] & !i[1821]) | ( l_47 [545] &  i[1821]);
assign l_46[273]    = ( l_47 [546] & !i[1821]) | ( l_47 [547] &  i[1821]);
assign l_46[274]    = ( l_47 [548] & !i[1821]) | ( l_47 [549] &  i[1821]);
assign l_46[275]    = ( l_47 [550] & !i[1821]) | ( l_47 [551] &  i[1821]);
assign l_46[276]    = ( l_47 [552] & !i[1821]) | ( l_47 [553] &  i[1821]);
assign l_46[277]    = ( l_47 [554] & !i[1821]) | ( l_47 [555] &  i[1821]);
assign l_46[278]    = ( l_47 [556] & !i[1821]) | ( l_47 [557] &  i[1821]);
assign l_46[279]    = ( l_47 [558] & !i[1821]) | ( l_47 [559] &  i[1821]);
assign l_46[280]    = ( l_47 [560] & !i[1821]) | ( l_47 [561] &  i[1821]);
assign l_46[281]    = ( l_47 [562] & !i[1821]) | ( l_47 [563] &  i[1821]);
assign l_46[282]    = ( l_47 [564] & !i[1821]) | ( l_47 [565] &  i[1821]);
assign l_46[283]    = ( l_47 [566] & !i[1821]) | ( l_47 [567] &  i[1821]);
assign l_46[284]    = ( l_47 [568] & !i[1821]) | ( l_47 [569] &  i[1821]);
assign l_46[285]    = ( l_47 [570] & !i[1821]) | ( l_47 [571] &  i[1821]);
assign l_46[286]    = ( l_47 [572] & !i[1821]) | ( l_47 [573] &  i[1821]);
assign l_46[287]    = ( l_47 [574] & !i[1821]) | ( l_47 [575] &  i[1821]);
assign l_46[288]    = ( l_47 [576] & !i[1821]) | ( l_47 [577] &  i[1821]);
assign l_46[289]    = ( l_47 [578] & !i[1821]) | ( l_47 [579] &  i[1821]);
assign l_46[290]    = ( l_47 [580] & !i[1821]) | ( l_47 [581] &  i[1821]);
assign l_46[291]    = ( l_47 [582] & !i[1821]) | ( l_47 [583] &  i[1821]);
assign l_46[292]    = ( l_47 [584] & !i[1821]) | ( l_47 [585] &  i[1821]);
assign l_46[293]    = ( l_47 [586] & !i[1821]) | ( l_47 [587] &  i[1821]);
assign l_46[294]    = ( l_47 [588] & !i[1821]) | ( l_47 [589] &  i[1821]);
assign l_46[295]    = ( l_47 [590] & !i[1821]) | ( l_47 [591] &  i[1821]);
assign l_46[296]    = ( l_47 [592] & !i[1821]) | ( l_47 [593] &  i[1821]);
assign l_46[297]    = ( l_47 [594] & !i[1821]) | ( l_47 [595] &  i[1821]);
assign l_46[298]    = ( l_47 [596] & !i[1821]) | ( l_47 [597] &  i[1821]);
assign l_46[299]    = ( l_47 [598] & !i[1821]) | ( l_47 [599] &  i[1821]);
assign l_46[300]    = ( l_47 [600] & !i[1821]) | ( l_47 [601] &  i[1821]);
assign l_46[301]    = ( l_47 [602] & !i[1821]) | ( l_47 [603] &  i[1821]);
assign l_46[302]    = ( l_47 [604] & !i[1821]) | ( l_47 [605] &  i[1821]);
assign l_46[303]    = ( l_47 [606] & !i[1821]) | ( l_47 [607] &  i[1821]);
assign l_46[304]    = ( l_47 [608] & !i[1821]) | ( l_47 [609] &  i[1821]);
assign l_46[305]    = ( l_47 [610] & !i[1821]) | ( l_47 [611] &  i[1821]);
assign l_46[306]    = ( l_47 [612] & !i[1821]) | ( l_47 [613] &  i[1821]);
assign l_46[307]    = ( l_47 [614] & !i[1821]) | ( l_47 [615] &  i[1821]);
assign l_46[308]    = ( l_47 [616] & !i[1821]) | ( l_47 [617] &  i[1821]);
assign l_46[309]    = ( l_47 [618] & !i[1821]) | ( l_47 [619] &  i[1821]);
assign l_46[310]    = ( l_47 [620] & !i[1821]) | ( l_47 [621] &  i[1821]);
assign l_46[311]    = ( l_47 [622] & !i[1821]) | ( l_47 [623] &  i[1821]);
assign l_46[312]    = ( l_47 [624] & !i[1821]) | ( l_47 [625] &  i[1821]);
assign l_46[313]    = ( l_47 [626] & !i[1821]) | ( l_47 [627] &  i[1821]);
assign l_46[314]    = ( l_47 [628] & !i[1821]) | ( l_47 [629] &  i[1821]);
assign l_46[315]    = ( l_47 [630] & !i[1821]) | ( l_47 [631] &  i[1821]);
assign l_46[316]    = ( l_47 [632] & !i[1821]) | ( l_47 [633] &  i[1821]);
assign l_46[317]    = ( l_47 [634] & !i[1821]) | ( l_47 [635] &  i[1821]);
assign l_46[318]    = ( l_47 [636] & !i[1821]) | ( l_47 [637] &  i[1821]);
assign l_46[319]    = ( l_47 [638] & !i[1821]) | ( l_47 [639] &  i[1821]);
assign l_46[320]    = ( l_47 [640] & !i[1821]) | ( l_47 [641] &  i[1821]);
assign l_46[321]    = ( l_47 [642] & !i[1821]) | ( l_47 [643] &  i[1821]);
assign l_46[322]    = ( l_47 [644] & !i[1821]) | ( l_47 [645] &  i[1821]);
assign l_46[323]    = ( l_47 [646] & !i[1821]) | ( l_47 [647] &  i[1821]);
assign l_46[324]    = ( l_47 [648] & !i[1821]) | ( l_47 [649] &  i[1821]);
assign l_46[325]    = ( l_47 [650] & !i[1821]) | ( l_47 [651] &  i[1821]);
assign l_46[326]    = ( l_47 [652] & !i[1821]) | ( l_47 [653] &  i[1821]);
assign l_46[327]    = ( l_47 [654] & !i[1821]) | ( l_47 [655] &  i[1821]);
assign l_46[328]    = ( l_47 [656]);
assign l_46[329]    = ( l_47 [657] & !i[1821]) | ( l_47 [658] &  i[1821]);
assign l_46[330]    = ( l_47 [659] & !i[1821]) | ( l_47 [660] &  i[1821]);
assign l_46[331]    = ( l_47 [661] & !i[1821]) | ( l_47 [662] &  i[1821]);
assign l_46[332]    = ( l_47 [663] & !i[1821]) | ( l_47 [664] &  i[1821]);
assign l_46[333]    = ( l_47 [665] & !i[1821]) | ( l_47 [666] &  i[1821]);
assign l_46[334]    = ( l_47 [667] & !i[1821]) | ( l_47 [668] &  i[1821]);
assign l_46[335]    = ( l_47 [669] & !i[1821]) | ( l_47 [670] &  i[1821]);
assign l_46[336]    = ( l_47 [671] & !i[1821]) | ( l_47 [672] &  i[1821]);
assign l_46[337]    = ( l_47 [673] & !i[1821]) | ( l_47 [674] &  i[1821]);
assign l_46[338]    = ( l_47 [675] & !i[1821]) | ( l_47 [676] &  i[1821]);
assign l_46[339]    = ( l_47 [677] & !i[1821]) | ( l_47 [678] &  i[1821]);
assign l_46[340]    = ( l_47 [679] & !i[1821]) | ( l_47 [680] &  i[1821]);
assign l_46[341]    = ( l_47 [681] & !i[1821]) | ( l_47 [682] &  i[1821]);
assign l_46[342]    = ( l_47 [683] & !i[1821]) | ( l_47 [684] &  i[1821]);
assign l_46[343]    = ( l_47 [685] & !i[1821]) | ( l_47 [686] &  i[1821]);
assign l_46[344]    = ( l_47 [687] & !i[1821]) | ( l_47 [688] &  i[1821]);
assign l_46[345]    = ( l_47 [689] & !i[1821]) | ( l_47 [690] &  i[1821]);
assign l_46[346]    = ( l_47 [691] & !i[1821]) | ( l_47 [692] &  i[1821]);
assign l_46[347]    = ( l_47 [693] & !i[1821]) | ( l_47 [694] &  i[1821]);
assign l_46[348]    = ( l_47 [695] & !i[1821]) | ( l_47 [696] &  i[1821]);
assign l_46[349]    = ( l_47 [697] & !i[1821]) | ( l_47 [698] &  i[1821]);
assign l_46[350]    = ( l_47 [699] & !i[1821]) | ( l_47 [700] &  i[1821]);
assign l_46[351]    = ( l_47 [701] & !i[1821]) | ( l_47 [702] &  i[1821]);
assign l_46[352]    = ( l_47 [703] & !i[1821]) | ( l_47 [704] &  i[1821]);
assign l_46[353]    = ( l_47 [705] & !i[1821]) | ( l_47 [706] &  i[1821]);
assign l_46[354]    = ( l_47 [707] & !i[1821]) | ( l_47 [708] &  i[1821]);
assign l_46[355]    = ( l_47 [709] & !i[1821]) | ( l_47 [710] &  i[1821]);
assign l_46[356]    = ( l_47 [711] & !i[1821]) | ( l_47 [712] &  i[1821]);
assign l_46[357]    = ( l_47 [713] & !i[1821]) | ( l_47 [714] &  i[1821]);
assign l_46[358]    = ( l_47 [715] & !i[1821]) | ( l_47 [716] &  i[1821]);
assign l_46[359]    = ( l_47 [717] & !i[1821]) | ( l_47 [718] &  i[1821]);
assign l_46[360]    = ( l_47 [719] & !i[1821]) | ( l_47 [720] &  i[1821]);
assign l_46[361]    = ( l_47 [721] & !i[1821]) | ( l_47 [722] &  i[1821]);
assign l_46[362]    = ( l_47 [723] & !i[1821]) | ( l_47 [724] &  i[1821]);
assign l_46[363]    = ( l_47 [725] & !i[1821]) | ( l_47 [726] &  i[1821]);
assign l_46[364]    = ( l_47 [727] & !i[1821]) | ( l_47 [728] &  i[1821]);
assign l_46[365]    = ( l_47 [729] & !i[1821]) | ( l_47 [730] &  i[1821]);
assign l_46[366]    = ( l_47 [731] & !i[1821]) | ( l_47 [732] &  i[1821]);
assign l_46[367]    = ( l_47 [733] & !i[1821]) | ( l_47 [734] &  i[1821]);
assign l_46[368]    = ( l_47 [735] & !i[1821]) | ( l_47 [736] &  i[1821]);
assign l_46[369]    = ( l_47 [737] & !i[1821]) | ( l_47 [738] &  i[1821]);
assign l_46[370]    = ( l_47 [739] & !i[1821]) | ( l_47 [740] &  i[1821]);
assign l_46[371]    = ( l_47 [741] & !i[1821]) | ( l_47 [742] &  i[1821]);
assign l_46[372]    = ( l_47 [743] & !i[1821]) | ( l_47 [744] &  i[1821]);
assign l_46[373]    = ( l_47 [745] & !i[1821]) | ( l_47 [746] &  i[1821]);
assign l_46[374]    = ( l_47 [747] & !i[1821]) | ( l_47 [748] &  i[1821]);
assign l_46[375]    = ( l_47 [749] & !i[1821]) | ( l_47 [750] &  i[1821]);
assign l_46[376]    = ( l_47 [751] & !i[1821]) | ( l_47 [752] &  i[1821]);
assign l_46[377]    = ( l_47 [753] & !i[1821]) | ( l_47 [754] &  i[1821]);
assign l_46[378]    = ( l_47 [755] & !i[1821]) | ( l_47 [756] &  i[1821]);
assign l_46[379]    = ( l_47 [757] & !i[1821]) | ( l_47 [758] &  i[1821]);
assign l_46[380]    = ( l_47 [759] & !i[1821]) | ( l_47 [760] &  i[1821]);
assign l_46[381]    = ( l_47 [761] & !i[1821]) | ( l_47 [762] &  i[1821]);
assign l_46[382]    = ( l_47 [763] & !i[1821]) | ( l_47 [764] &  i[1821]);
assign l_46[383]    = ( l_47 [765] & !i[1821]) | ( l_47 [766] &  i[1821]);
assign l_46[384]    = ( l_47 [767] & !i[1821]) | ( l_47 [768] &  i[1821]);
assign l_46[385]    = ( l_47 [769] & !i[1821]) | ( l_47 [770] &  i[1821]);
assign l_46[386]    = ( l_47 [771] & !i[1821]) | ( l_47 [772] &  i[1821]);
assign l_46[387]    = ( l_47 [773] & !i[1821]) | ( l_47 [774] &  i[1821]);
assign l_46[388]    = ( l_47 [775] & !i[1821]) | ( l_47 [776] &  i[1821]);
assign l_46[389]    = ( l_47 [777] & !i[1821]) | ( l_47 [778] &  i[1821]);
assign l_46[390]    = ( l_47 [779] & !i[1821]) | ( l_47 [780] &  i[1821]);
assign l_46[391]    = ( l_47 [781] & !i[1821]) | ( l_47 [782] &  i[1821]);
assign l_46[392]    = ( l_47 [783] & !i[1821]) | ( l_47 [784] &  i[1821]);
assign l_46[393]    = ( l_47 [785] & !i[1821]) | ( l_47 [786] &  i[1821]);
assign l_46[394]    = ( l_47 [787] & !i[1821]) | ( l_47 [788] &  i[1821]);
assign l_46[395]    = ( l_47 [789] & !i[1821]) | ( l_47 [790] &  i[1821]);
assign l_46[396]    = ( l_47 [791] & !i[1821]) | ( l_47 [792] &  i[1821]);
assign l_46[397]    = ( l_47 [793] & !i[1821]) | ( l_47 [794] &  i[1821]);
assign l_46[398]    = ( l_47 [795] & !i[1821]) | ( l_47 [796] &  i[1821]);
assign l_46[399]    = ( l_47 [797] & !i[1821]) | ( l_47 [798] &  i[1821]);
assign l_46[400]    = ( l_47 [799] & !i[1821]) | ( l_47 [800] &  i[1821]);
assign l_46[401]    = ( l_47 [801] & !i[1821]) | ( l_47 [802] &  i[1821]);
assign l_46[402]    = ( l_47 [803] & !i[1821]) | ( l_47 [804] &  i[1821]);
assign l_46[403]    = ( l_47 [805] & !i[1821]) | ( l_47 [806] &  i[1821]);
assign l_46[404]    = ( l_47 [807] & !i[1821]) | ( l_47 [808] &  i[1821]);
assign l_46[405]    = ( l_47 [809] & !i[1821]) | ( l_47 [810] &  i[1821]);
assign l_46[406]    = ( l_47 [811] & !i[1821]) | ( l_47 [812] &  i[1821]);
assign l_46[407]    = ( l_47 [813] & !i[1821]) | ( l_47 [814] &  i[1821]);
assign l_46[408]    = ( l_47 [815] & !i[1821]) | ( l_47 [816] &  i[1821]);
assign l_46[409]    = ( l_47 [817] & !i[1821]) | ( l_47 [818] &  i[1821]);
assign l_46[410]    = ( l_47 [819] & !i[1821]) | ( l_47 [820] &  i[1821]);
assign l_46[411]    = ( l_47 [821] & !i[1821]) | ( l_47 [822] &  i[1821]);
assign l_46[412]    = ( l_47 [823] & !i[1821]) | ( l_47 [824] &  i[1821]);
assign l_46[413]    = ( l_47 [825] & !i[1821]) | ( l_47 [826] &  i[1821]);
assign l_46[414]    = ( l_47 [827] & !i[1821]) | ( l_47 [828] &  i[1821]);
assign l_46[415]    = ( l_47 [829] & !i[1821]) | ( l_47 [830] &  i[1821]);
assign l_46[416]    = ( l_47 [831] & !i[1821]) | ( l_47 [832] &  i[1821]);
assign l_46[417]    = ( l_47 [833] & !i[1821]) | ( l_47 [834] &  i[1821]);
assign l_46[418]    = ( l_47 [835] & !i[1821]) | ( l_47 [836] &  i[1821]);
assign l_46[419]    = ( l_47 [837] & !i[1821]) | ( l_47 [838] &  i[1821]);
assign l_46[420]    = ( l_47 [839] & !i[1821]) | ( l_47 [840] &  i[1821]);
assign l_46[421]    = ( l_47 [841] & !i[1821]) | ( l_47 [842] &  i[1821]);
assign l_46[422]    = ( l_47 [843] & !i[1821]) | ( l_47 [844] &  i[1821]);
assign l_46[423]    = ( l_47 [845] & !i[1821]) | ( l_47 [846] &  i[1821]);
assign l_46[424]    = ( l_47 [847] & !i[1821]) | ( l_47 [848] &  i[1821]);
assign l_46[425]    = ( l_47 [849] & !i[1821]) | ( l_47 [850] &  i[1821]);
assign l_46[426]    = ( l_47 [851] & !i[1821]) | ( l_47 [852] &  i[1821]);
assign l_46[427]    = ( l_47 [853] & !i[1821]) | ( l_47 [854] &  i[1821]);
assign l_46[428]    = ( l_47 [855] & !i[1821]) | ( l_47 [856] &  i[1821]);
assign l_46[429]    = ( l_47 [857] & !i[1821]) | ( l_47 [858] &  i[1821]);
assign l_46[430]    = ( l_47 [859] & !i[1821]) | ( l_47 [860] &  i[1821]);
assign l_46[431]    = ( l_47 [861] & !i[1821]) | ( l_47 [862] &  i[1821]);
assign l_46[432]    = ( l_47 [863] & !i[1821]) | ( l_47 [864] &  i[1821]);
assign l_46[433]    = ( l_47 [865] & !i[1821]) | ( l_47 [866] &  i[1821]);
assign l_46[434]    = ( l_47 [867] & !i[1821]) | ( l_47 [868] &  i[1821]);
assign l_46[435]    = ( l_47 [869] & !i[1821]) | ( l_47 [870] &  i[1821]);
assign l_46[436]    = ( l_47 [871] & !i[1821]) | ( l_47 [872] &  i[1821]);
assign l_46[437]    = ( l_47 [873] & !i[1821]) | ( l_47 [874] &  i[1821]);
assign l_46[438]    = ( l_47 [875] & !i[1821]) | ( l_47 [876] &  i[1821]);
assign l_46[439]    = ( l_47 [877] & !i[1821]) | ( l_47 [878] &  i[1821]);
assign l_46[440]    = ( l_47 [879] & !i[1821]) | ( l_47 [880] &  i[1821]);
assign l_46[441]    = ( l_47 [881] & !i[1821]) | ( l_47 [882] &  i[1821]);
assign l_46[442]    = ( l_47 [883] & !i[1821]) | ( l_47 [884] &  i[1821]);
assign l_46[443]    = ( l_47 [885] & !i[1821]) | ( l_47 [886] &  i[1821]);
assign l_46[444]    = ( l_47 [887] & !i[1821]) | ( l_47 [888] &  i[1821]);
assign l_46[445]    = ( l_47 [889] & !i[1821]) | ( l_47 [890] &  i[1821]);
assign l_46[446]    = ( l_47 [891] & !i[1821]) | ( l_47 [892] &  i[1821]);
assign l_46[447]    = ( l_47 [893] & !i[1821]) | ( l_47 [894] &  i[1821]);
assign l_46[448]    = ( l_47 [895] & !i[1821]) | ( l_47 [896] &  i[1821]);
assign l_46[449]    = ( l_47 [897] & !i[1821]) | ( l_47 [898] &  i[1821]);
assign l_46[450]    = ( l_47 [899] & !i[1821]) | ( l_47 [900] &  i[1821]);
assign l_46[451]    = ( l_47 [901] & !i[1821]) | ( l_47 [902] &  i[1821]);
assign l_46[452]    = ( l_47 [903] & !i[1821]) | ( l_47 [904] &  i[1821]);
assign l_46[453]    = ( l_47 [905] & !i[1821]) | ( l_47 [906] &  i[1821]);
assign l_46[454]    = ( l_47 [907] & !i[1821]) | ( l_47 [908] &  i[1821]);
assign l_46[455]    = ( l_47 [909] & !i[1821]) | ( l_47 [910] &  i[1821]);
assign l_46[456]    = ( l_47 [911] & !i[1821]) | ( l_47 [912] &  i[1821]);
assign l_46[457]    = ( l_47 [913] & !i[1821]) | ( l_47 [914] &  i[1821]);
assign l_46[458]    = ( l_47 [915] & !i[1821]) | ( l_47 [916] &  i[1821]);
assign l_46[459]    = ( l_47 [917] & !i[1821]) | ( l_47 [918] &  i[1821]);
assign l_46[460]    = ( l_47 [919] & !i[1821]) | ( l_47 [920] &  i[1821]);
assign l_46[461]    = ( l_47 [921] & !i[1821]) | ( l_47 [922] &  i[1821]);
assign l_46[462]    = ( l_47 [923] & !i[1821]) | ( l_47 [924] &  i[1821]);
assign l_46[463]    = ( l_47 [925] & !i[1821]) | ( l_47 [926] &  i[1821]);
assign l_46[464]    = ( l_47 [927] & !i[1821]) | ( l_47 [928] &  i[1821]);
assign l_46[465]    = ( l_47 [929] & !i[1821]) | ( l_47 [930] &  i[1821]);
assign l_46[466]    = ( l_47 [931] & !i[1821]) | ( l_47 [932] &  i[1821]);
assign l_46[467]    = ( l_47 [933] & !i[1821]) | ( l_47 [934] &  i[1821]);
assign l_46[468]    = ( l_47 [935] & !i[1821]) | ( l_47 [936] &  i[1821]);
assign l_46[469]    = ( l_47 [937] & !i[1821]) | ( l_47 [938] &  i[1821]);
assign l_46[470]    = ( l_47 [939] & !i[1821]) | ( l_47 [940] &  i[1821]);
assign l_46[471]    = ( l_47 [941] & !i[1821]) | ( l_47 [942] &  i[1821]);
assign l_46[472]    = ( l_47 [943] & !i[1821]) | ( l_47 [944] &  i[1821]);
assign l_46[473]    = ( l_47 [945] & !i[1821]) | ( l_47 [946] &  i[1821]);
assign l_46[474]    = ( l_47 [947] & !i[1821]) | ( l_47 [948] &  i[1821]);
assign l_46[475]    = ( l_47 [949] & !i[1821]) | ( l_47 [950] &  i[1821]);
assign l_46[476]    = ( l_47 [951] & !i[1821]) | ( l_47 [952] &  i[1821]);
assign l_46[477]    = ( l_47 [953] & !i[1821]) | ( l_47 [954] &  i[1821]);
assign l_46[478]    = ( l_47 [955] & !i[1821]) | ( l_47 [956] &  i[1821]);
assign l_46[479]    = ( l_47 [957] & !i[1821]) | ( l_47 [958] &  i[1821]);
assign l_46[480]    = ( l_47 [959] & !i[1821]) | ( l_47 [960] &  i[1821]);
assign l_46[481]    = ( l_47 [961] & !i[1821]) | ( l_47 [962] &  i[1821]);
assign l_46[482]    = ( l_47 [963] & !i[1821]) | ( l_47 [964] &  i[1821]);
assign l_46[483]    = ( l_47 [965] & !i[1821]) | ( l_47 [966] &  i[1821]);
assign l_46[484]    = ( l_47 [967] & !i[1821]) | ( l_47 [968] &  i[1821]);
assign l_46[485]    = ( l_47 [969] & !i[1821]) | ( l_47 [970] &  i[1821]);
assign l_46[486]    = ( l_47 [971] & !i[1821]) | ( l_47 [972] &  i[1821]);
assign l_46[487]    = ( l_47 [973] & !i[1821]) | ( l_47 [974] &  i[1821]);
assign l_46[488]    = ( l_47 [975] & !i[1821]) | ( l_47 [976] &  i[1821]);
assign l_46[489]    = ( l_47 [977] & !i[1821]) | ( l_47 [978] &  i[1821]);
assign l_46[490]    = ( l_47 [979] & !i[1821]) | ( l_47 [980] &  i[1821]);
assign l_46[491]    = ( l_47 [981] & !i[1821]) | ( l_47 [982] &  i[1821]);
assign l_46[492]    = ( l_47 [983] & !i[1821]) | ( l_47 [984] &  i[1821]);
assign l_46[493]    = ( l_47 [985] & !i[1821]) | ( l_47 [986] &  i[1821]);
assign l_46[494]    = ( l_47 [987] & !i[1821]) | ( l_47 [988] &  i[1821]);
assign l_46[495]    = ( l_47 [989] & !i[1821]) | ( l_47 [990] &  i[1821]);
assign l_46[496]    = ( l_47 [991] & !i[1821]) | ( l_47 [992] &  i[1821]);
assign l_46[497]    = ( l_47 [993] & !i[1821]) | ( l_47 [994] &  i[1821]);
assign l_46[498]    = ( l_47 [995] & !i[1821]) | ( l_47 [996] &  i[1821]);
assign l_46[499]    = ( l_47 [997] & !i[1821]) | ( l_47 [998] &  i[1821]);
assign l_46[500]    = ( l_47 [999] & !i[1821]) | ( l_47 [1000] &  i[1821]);
assign l_46[501]    = ( l_47 [1001] & !i[1821]) | ( l_47 [1002] &  i[1821]);
assign l_46[502]    = ( l_47 [1003] & !i[1821]) | ( l_47 [1004] &  i[1821]);
assign l_46[503]    = ( l_47 [1005] & !i[1821]) | ( l_47 [1006] &  i[1821]);
assign l_46[504]    = ( l_47 [1007] & !i[1821]) | ( l_47 [1008] &  i[1821]);
assign l_46[505]    = ( l_47 [1009] & !i[1821]) | ( l_47 [1010] &  i[1821]);
assign l_46[506]    = ( l_47 [1011] & !i[1821]) | ( l_47 [1012] &  i[1821]);
assign l_46[507]    = ( l_47 [1013] & !i[1821]) | ( l_47 [1014] &  i[1821]);
assign l_46[508]    = ( l_47 [1015] & !i[1821]) | ( l_47 [1016] &  i[1821]);
assign l_46[509]    = ( l_47 [1017] & !i[1821]) | ( l_47 [1018] &  i[1821]);
assign l_46[510]    = ( l_47 [1019] & !i[1821]) | ( l_47 [1020] &  i[1821]);
assign l_46[511]    = ( l_47 [1021] & !i[1821]) | ( l_47 [1022] &  i[1821]);
assign l_46[512]    = ( l_47 [1023] & !i[1821]) | ( l_47 [1024] &  i[1821]);
assign l_46[513]    = ( l_47 [1025] & !i[1821]) | ( l_47 [1026] &  i[1821]);
assign l_46[514]    = ( l_47 [1027] & !i[1821]) | ( l_47 [1028] &  i[1821]);
assign l_46[515]    = ( l_47 [1029] & !i[1821]) | ( l_47 [1030] &  i[1821]);
assign l_46[516]    = ( l_47 [1031] & !i[1821]) | ( l_47 [1032] &  i[1821]);
assign l_46[517]    = ( l_47 [1033] & !i[1821]) | ( l_47 [1034] &  i[1821]);
assign l_46[518]    = ( l_47 [1035] & !i[1821]) | ( l_47 [1036] &  i[1821]);
assign l_46[519]    = ( l_47 [1037] & !i[1821]) | ( l_47 [1038] &  i[1821]);
assign l_46[520]    = ( l_47 [1039] & !i[1821]) | ( l_47 [1040] &  i[1821]);
assign l_46[521]    = ( l_47 [1041] & !i[1821]) | ( l_47 [1042] &  i[1821]);
assign l_46[522]    = ( l_47 [1043] & !i[1821]) | ( l_47 [1044] &  i[1821]);
assign l_46[523]    = ( l_47 [1045] & !i[1821]) | ( l_47 [1046] &  i[1821]);
assign l_46[524]    = ( l_47 [1047] & !i[1821]) | ( l_47 [1048] &  i[1821]);
assign l_46[525]    = ( l_47 [1049] & !i[1821]) | ( l_47 [1050] &  i[1821]);
assign l_46[526]    = ( l_47 [1051] & !i[1821]) | ( l_47 [1052] &  i[1821]);
assign l_46[527]    = ( l_47 [1053] & !i[1821]) | ( l_47 [1054] &  i[1821]);
assign l_46[528]    = ( l_47 [1055] & !i[1821]) | ( l_47 [1056] &  i[1821]);
assign l_46[529]    = ( l_47 [1057]);
assign l_46[530]    = ( l_47 [1058]);
assign l_46[531]    = ( l_47 [1059]);
assign l_46[532]    =  i[1821];
assign l_46[533]    = ( l_47 [1060]);
assign l_46[534]    = ( l_47 [1061]);
assign l_46[535]    = ( l_47 [1062]);
assign l_46[536]    = ( l_47 [1063]);
assign l_47[0]    = ( l_48 [0] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[1]    = ( l_48 [2] & !i[1699]) | ( l_48 [0] &  i[1699]);
assign l_47[2]    = ( l_48 [3] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[3]    = ( l_48 [2] & !i[1699]) | ( l_48 [3] &  i[1699]);
assign l_47[4]    = ( l_48 [4] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[5]    = ( l_48 [2] & !i[1699]) | ( l_48 [4] &  i[1699]);
assign l_47[6]    = ( l_48 [5] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[7]    = ( l_48 [2] & !i[1699]) | ( l_48 [5] &  i[1699]);
assign l_47[8]    = ( l_48 [6] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[9]    = ( l_48 [2] & !i[1699]) | ( l_48 [6] &  i[1699]);
assign l_47[10]    = ( l_48 [7] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[11]    = ( l_48 [2] & !i[1699]) | ( l_48 [7] &  i[1699]);
assign l_47[12]    = ( l_48 [8] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[13]    = ( l_48 [2] & !i[1699]) | ( l_48 [8] &  i[1699]);
assign l_47[14]    = ( l_48 [9] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[15]    = ( l_48 [2] & !i[1699]) | ( l_48 [9] &  i[1699]);
assign l_47[16]    = ( l_48 [10] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[17]    = ( l_48 [2] & !i[1699]) | ( l_48 [10] &  i[1699]);
assign l_47[18]    = ( l_48 [11] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[19]    = ( l_48 [2] & !i[1699]) | ( l_48 [11] &  i[1699]);
assign l_47[20]    = ( l_48 [12] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[21]    = ( l_48 [2] & !i[1699]) | ( l_48 [12] &  i[1699]);
assign l_47[22]    = ( l_48 [13] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[23]    = ( l_48 [2] & !i[1699]) | ( l_48 [13] &  i[1699]);
assign l_47[24]    = ( l_48 [14] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[25]    = ( l_48 [2] & !i[1699]) | ( l_48 [14] &  i[1699]);
assign l_47[26]    = ( l_48 [15] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[27]    = ( l_48 [2] & !i[1699]) | ( l_48 [15] &  i[1699]);
assign l_47[28]    = ( l_48 [16] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[29]    = ( l_48 [2] & !i[1699]) | ( l_48 [16] &  i[1699]);
assign l_47[30]    = ( l_48 [17] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[31]    = ( l_48 [2] & !i[1699]) | ( l_48 [17] &  i[1699]);
assign l_47[32]    = ( l_48 [18] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[33]    = ( l_48 [19] & !i[1699]) | ( l_48 [18] &  i[1699]);
assign l_47[34]    = ( l_48 [20] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[35]    = ( l_48 [19] & !i[1699]) | ( l_48 [20] &  i[1699]);
assign l_47[36]    = ( l_48 [21] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[37]    = ( l_48 [19] & !i[1699]) | ( l_48 [21] &  i[1699]);
assign l_47[38]    = ( l_48 [22] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[39]    = ( l_48 [19] & !i[1699]) | ( l_48 [22] &  i[1699]);
assign l_47[40]    = ( l_48 [23] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[41]    = ( l_48 [19] & !i[1699]) | ( l_48 [23] &  i[1699]);
assign l_47[42]    = ( l_48 [24] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[43]    = ( l_48 [19] & !i[1699]) | ( l_48 [24] &  i[1699]);
assign l_47[44]    = ( l_48 [25] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[45]    = ( l_48 [19] & !i[1699]) | ( l_48 [25] &  i[1699]);
assign l_47[46]    = ( l_48 [26] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[47]    = ( l_48 [19] & !i[1699]) | ( l_48 [26] &  i[1699]);
assign l_47[48]    = ( l_48 [27] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[49]    = ( l_48 [19] & !i[1699]) | ( l_48 [27] &  i[1699]);
assign l_47[50]    = ( l_48 [28] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[51]    = ( l_48 [19] & !i[1699]) | ( l_48 [28] &  i[1699]);
assign l_47[52]    = ( l_48 [29] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[53]    = ( l_48 [19] & !i[1699]) | ( l_48 [29] &  i[1699]);
assign l_47[54]    = ( l_48 [30] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[55]    = ( l_48 [19] & !i[1699]) | ( l_48 [30] &  i[1699]);
assign l_47[56]    = ( l_48 [31] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[57]    = ( l_48 [19] & !i[1699]) | ( l_48 [31] &  i[1699]);
assign l_47[58]    = ( l_48 [32] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[59]    = ( l_48 [19] & !i[1699]) | ( l_48 [32] &  i[1699]);
assign l_47[60]    = ( l_48 [33] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[61]    = ( l_48 [19] & !i[1699]) | ( l_48 [33] &  i[1699]);
assign l_47[62]    = ( l_48 [34] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[63]    = ( l_48 [19] & !i[1699]) | ( l_48 [34] &  i[1699]);
assign l_47[64]    = ( l_48 [35] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[65]    = ( l_48 [36] & !i[1699]) | ( l_48 [35] &  i[1699]);
assign l_47[66]    = ( l_48 [37] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[67]    = ( l_48 [36] & !i[1699]) | ( l_48 [37] &  i[1699]);
assign l_47[68]    = ( l_48 [38] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[69]    = ( l_48 [36] & !i[1699]) | ( l_48 [38] &  i[1699]);
assign l_47[70]    = ( l_48 [39] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[71]    = ( l_48 [36] & !i[1699]) | ( l_48 [39] &  i[1699]);
assign l_47[72]    = ( l_48 [40] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[73]    = ( l_48 [36] & !i[1699]) | ( l_48 [40] &  i[1699]);
assign l_47[74]    = ( l_48 [41] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[75]    = ( l_48 [36] & !i[1699]) | ( l_48 [41] &  i[1699]);
assign l_47[76]    = ( l_48 [42] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[77]    = ( l_48 [36] & !i[1699]) | ( l_48 [42] &  i[1699]);
assign l_47[78]    = ( l_48 [43] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[79]    = ( l_48 [36] & !i[1699]) | ( l_48 [43] &  i[1699]);
assign l_47[80]    = ( l_48 [44] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[81]    = ( l_48 [36] & !i[1699]) | ( l_48 [44] &  i[1699]);
assign l_47[82]    = ( l_48 [45] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[83]    = ( l_48 [36] & !i[1699]) | ( l_48 [45] &  i[1699]);
assign l_47[84]    = ( l_48 [46] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[85]    = ( l_48 [36] & !i[1699]) | ( l_48 [46] &  i[1699]);
assign l_47[86]    = ( l_48 [47] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[87]    = ( l_48 [36] & !i[1699]) | ( l_48 [47] &  i[1699]);
assign l_47[88]    = ( l_48 [48] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[89]    = ( l_48 [36] & !i[1699]) | ( l_48 [48] &  i[1699]);
assign l_47[90]    = ( l_48 [49] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[91]    = ( l_48 [36] & !i[1699]) | ( l_48 [49] &  i[1699]);
assign l_47[92]    = ( l_48 [50] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[93]    = ( l_48 [36] & !i[1699]) | ( l_48 [50] &  i[1699]);
assign l_47[94]    = ( l_48 [51] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[95]    = ( l_48 [36] & !i[1699]) | ( l_48 [51] &  i[1699]);
assign l_47[96]    = ( l_48 [52] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[97]    = ( l_48 [52] &  i[1699]);
assign l_47[98]    = ( l_48 [53] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[99]    = ( l_48 [53] &  i[1699]);
assign l_47[100]    = ( l_48 [54] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[101]    = ( l_48 [54] &  i[1699]);
assign l_47[102]    = ( l_48 [55] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[103]    = ( l_48 [55] &  i[1699]);
assign l_47[104]    = ( l_48 [56] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[105]    = ( l_48 [56] &  i[1699]);
assign l_47[106]    = ( l_48 [57] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[107]    = ( l_48 [57] &  i[1699]);
assign l_47[108]    = ( l_48 [58] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[109]    = ( l_48 [58] &  i[1699]);
assign l_47[110]    = ( l_48 [59] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[111]    = ( l_48 [59] &  i[1699]);
assign l_47[112]    = ( l_48 [60] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[113]    = ( l_48 [60] &  i[1699]);
assign l_47[114]    = ( l_48 [61] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[115]    = ( l_48 [61] &  i[1699]);
assign l_47[116]    = ( l_48 [62] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[117]    = ( l_48 [62] &  i[1699]);
assign l_47[118]    = ( l_48 [63] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[119]    = ( l_48 [63] &  i[1699]);
assign l_47[120]    = ( l_48 [64] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[121]    = ( l_48 [64] &  i[1699]);
assign l_47[122]    = ( l_48 [65] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[123]    = ( l_48 [65] &  i[1699]);
assign l_47[124]    = ( l_48 [66] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[125]    = ( l_48 [66] &  i[1699]);
assign l_47[126]    = ( l_48 [67] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[127]    = ( l_48 [67] &  i[1699]);
assign l_47[128]    = ( l_48 [68] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[129]    = ( l_48 [2] & !i[1699]) | ( l_48 [68] &  i[1699]);
assign l_47[130]    = ( l_48 [69] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[131]    = ( l_48 [2] & !i[1699]) | ( l_48 [69] &  i[1699]);
assign l_47[132]    = ( l_48 [70] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[133]    = ( l_48 [2] & !i[1699]) | ( l_48 [70] &  i[1699]);
assign l_47[134]    = ( l_48 [71] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[135]    = ( l_48 [2] & !i[1699]) | ( l_48 [71] &  i[1699]);
assign l_47[136]    = ( l_48 [72] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[137]    = ( l_48 [2] & !i[1699]) | ( l_48 [72] &  i[1699]);
assign l_47[138]    = ( l_48 [73] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[139]    = ( l_48 [2] & !i[1699]) | ( l_48 [73] &  i[1699]);
assign l_47[140]    = ( l_48 [74] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[141]    = ( l_48 [2] & !i[1699]) | ( l_48 [74] &  i[1699]);
assign l_47[142]    = ( l_48 [75] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[143]    = ( l_48 [2] & !i[1699]) | ( l_48 [75] &  i[1699]);
assign l_47[144]    = ( l_48 [76] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[145]    = ( l_48 [2] & !i[1699]) | ( l_48 [76] &  i[1699]);
assign l_47[146]    = ( l_48 [77] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[147]    = ( l_48 [2] & !i[1699]) | ( l_48 [77] &  i[1699]);
assign l_47[148]    = ( l_48 [78] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[149]    = ( l_48 [2] & !i[1699]) | ( l_48 [78] &  i[1699]);
assign l_47[150]    = ( l_48 [79] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[151]    = ( l_48 [2] & !i[1699]) | ( l_48 [79] &  i[1699]);
assign l_47[152]    = ( l_48 [80] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[153]    = ( l_48 [2] & !i[1699]) | ( l_48 [80] &  i[1699]);
assign l_47[154]    = ( l_48 [81] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[155]    = ( l_48 [2] & !i[1699]) | ( l_48 [81] &  i[1699]);
assign l_47[156]    = ( l_48 [82] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[157]    = ( l_48 [2] & !i[1699]) | ( l_48 [82] &  i[1699]);
assign l_47[158]    = ( l_48 [83] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[159]    = ( l_48 [2] & !i[1699]) | ( l_48 [83] &  i[1699]);
assign l_47[160]    = ( l_48 [84] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[161]    = ( l_48 [19] & !i[1699]) | ( l_48 [84] &  i[1699]);
assign l_47[162]    = ( l_48 [85] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[163]    = ( l_48 [19] & !i[1699]) | ( l_48 [85] &  i[1699]);
assign l_47[164]    = ( l_48 [86] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[165]    = ( l_48 [19] & !i[1699]) | ( l_48 [86] &  i[1699]);
assign l_47[166]    = ( l_48 [87] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[167]    = ( l_48 [19] & !i[1699]) | ( l_48 [87] &  i[1699]);
assign l_47[168]    = ( l_48 [88] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[169]    = ( l_48 [19] & !i[1699]) | ( l_48 [88] &  i[1699]);
assign l_47[170]    = ( l_48 [89] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[171]    = ( l_48 [19] & !i[1699]) | ( l_48 [89] &  i[1699]);
assign l_47[172]    = ( l_48 [90] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[173]    = ( l_48 [19] & !i[1699]) | ( l_48 [90] &  i[1699]);
assign l_47[174]    = ( l_48 [91] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[175]    = ( l_48 [19] & !i[1699]) | ( l_48 [91] &  i[1699]);
assign l_47[176]    = ( l_48 [92] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[177]    = ( l_48 [19] & !i[1699]) | ( l_48 [92] &  i[1699]);
assign l_47[178]    = ( l_48 [93] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[179]    = ( l_48 [19] & !i[1699]) | ( l_48 [93] &  i[1699]);
assign l_47[180]    = ( l_48 [94] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[181]    = ( l_48 [19] & !i[1699]) | ( l_48 [94] &  i[1699]);
assign l_47[182]    = ( l_48 [95] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[183]    = ( l_48 [19] & !i[1699]) | ( l_48 [95] &  i[1699]);
assign l_47[184]    = ( l_48 [96] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[185]    = ( l_48 [19] & !i[1699]) | ( l_48 [96] &  i[1699]);
assign l_47[186]    = ( l_48 [97] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[187]    = ( l_48 [19] & !i[1699]) | ( l_48 [97] &  i[1699]);
assign l_47[188]    = ( l_48 [98] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[189]    = ( l_48 [19] & !i[1699]) | ( l_48 [98] &  i[1699]);
assign l_47[190]    = ( l_48 [99] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[191]    = ( l_48 [19] & !i[1699]) | ( l_48 [99] &  i[1699]);
assign l_47[192]    = ( l_48 [100] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[193]    = ( l_48 [36] & !i[1699]) | ( l_48 [100] &  i[1699]);
assign l_47[194]    = ( l_48 [101] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[195]    = ( l_48 [36] & !i[1699]) | ( l_48 [101] &  i[1699]);
assign l_47[196]    = ( l_48 [102] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[197]    = ( l_48 [36] & !i[1699]) | ( l_48 [102] &  i[1699]);
assign l_47[198]    = ( l_48 [103] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[199]    = ( l_48 [36] & !i[1699]) | ( l_48 [103] &  i[1699]);
assign l_47[200]    = ( l_48 [104] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[201]    = ( l_48 [36] & !i[1699]) | ( l_48 [104] &  i[1699]);
assign l_47[202]    = ( l_48 [105] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[203]    = ( l_48 [36] & !i[1699]) | ( l_48 [105] &  i[1699]);
assign l_47[204]    = ( l_48 [106] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[205]    = ( l_48 [36] & !i[1699]) | ( l_48 [106] &  i[1699]);
assign l_47[206]    = ( l_48 [107] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[207]    = ( l_48 [36] & !i[1699]) | ( l_48 [107] &  i[1699]);
assign l_47[208]    = ( l_48 [108] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[209]    = ( l_48 [36] & !i[1699]) | ( l_48 [108] &  i[1699]);
assign l_47[210]    = ( l_48 [109] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[211]    = ( l_48 [36] & !i[1699]) | ( l_48 [109] &  i[1699]);
assign l_47[212]    = ( l_48 [110] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[213]    = ( l_48 [36] & !i[1699]) | ( l_48 [110] &  i[1699]);
assign l_47[214]    = ( l_48 [111] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[215]    = ( l_48 [36] & !i[1699]) | ( l_48 [111] &  i[1699]);
assign l_47[216]    = ( l_48 [112] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[217]    = ( l_48 [36] & !i[1699]) | ( l_48 [112] &  i[1699]);
assign l_47[218]    = ( l_48 [113] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[219]    = ( l_48 [36] & !i[1699]) | ( l_48 [113] &  i[1699]);
assign l_47[220]    = ( l_48 [114] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[221]    = ( l_48 [36] & !i[1699]) | ( l_48 [114] &  i[1699]);
assign l_47[222]    = ( l_48 [115] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[223]    = ( l_48 [36] & !i[1699]) | ( l_48 [115] &  i[1699]);
assign l_47[224]    = ( l_48 [116] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[225]    = ( l_48 [116] &  i[1699]);
assign l_47[226]    = ( l_48 [117] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[227]    = ( l_48 [117] &  i[1699]);
assign l_47[228]    = ( l_48 [118] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[229]    = ( l_48 [118] &  i[1699]);
assign l_47[230]    = ( l_48 [119] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[231]    = ( l_48 [119] &  i[1699]);
assign l_47[232]    = ( l_48 [120] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[233]    = ( l_48 [120] &  i[1699]);
assign l_47[234]    = ( l_48 [121] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[235]    = ( l_48 [121] &  i[1699]);
assign l_47[236]    = ( l_48 [122] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[237]    = ( l_48 [122] &  i[1699]);
assign l_47[238]    = ( l_48 [123] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[239]    = ( l_48 [123] &  i[1699]);
assign l_47[240]    = ( l_48 [124] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[241]    = ( l_48 [124] &  i[1699]);
assign l_47[242]    = ( l_48 [125] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[243]    = ( l_48 [125] &  i[1699]);
assign l_47[244]    = ( l_48 [126] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[245]    = ( l_48 [126] &  i[1699]);
assign l_47[246]    = ( l_48 [127] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[247]    = ( l_48 [127] &  i[1699]);
assign l_47[248]    = ( l_48 [128] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[249]    = ( l_48 [128] &  i[1699]);
assign l_47[250]    = ( l_48 [129] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[251]    = ( l_48 [129] &  i[1699]);
assign l_47[252]    = ( l_48 [130] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[253]    = ( l_48 [130] &  i[1699]);
assign l_47[254]    = ( l_48 [131] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[255]    = ( l_48 [131] &  i[1699]);
assign l_47[256]    = ( l_48 [132] & !i[1699]) | (      i[1699]);
assign l_47[257]    = ( l_48 [133] & !i[1699]) | ( l_48 [132] &  i[1699]);
assign l_47[258]    = ( l_48 [134] & !i[1699]) | (      i[1699]);
assign l_47[259]    = ( l_48 [133] & !i[1699]) | ( l_48 [134] &  i[1699]);
assign l_47[260]    = ( l_48 [135] & !i[1699]) | (      i[1699]);
assign l_47[261]    = ( l_48 [133] & !i[1699]) | ( l_48 [135] &  i[1699]);
assign l_47[262]    = ( l_48 [136] & !i[1699]) | (      i[1699]);
assign l_47[263]    = ( l_48 [133] & !i[1699]) | ( l_48 [136] &  i[1699]);
assign l_47[264]    = ( l_48 [137] & !i[1699]) | (      i[1699]);
assign l_47[265]    = ( l_48 [133] & !i[1699]) | ( l_48 [137] &  i[1699]);
assign l_47[266]    = ( l_48 [138] & !i[1699]) | (      i[1699]);
assign l_47[267]    = ( l_48 [133] & !i[1699]) | ( l_48 [138] &  i[1699]);
assign l_47[268]    = ( l_48 [139] & !i[1699]) | (      i[1699]);
assign l_47[269]    = ( l_48 [133] & !i[1699]) | ( l_48 [139] &  i[1699]);
assign l_47[270]    = ( l_48 [140] & !i[1699]) | (      i[1699]);
assign l_47[271]    = ( l_48 [133] & !i[1699]) | ( l_48 [140] &  i[1699]);
assign l_47[272]    = ( l_48 [141] & !i[1699]) | (      i[1699]);
assign l_47[273]    = ( l_48 [133] & !i[1699]) | ( l_48 [141] &  i[1699]);
assign l_47[274]    = ( l_48 [142] & !i[1699]) | (      i[1699]);
assign l_47[275]    = ( l_48 [133] & !i[1699]) | ( l_48 [142] &  i[1699]);
assign l_47[276]    = ( l_48 [143] & !i[1699]) | (      i[1699]);
assign l_47[277]    = ( l_48 [133] & !i[1699]) | ( l_48 [143] &  i[1699]);
assign l_47[278]    = ( l_48 [144] & !i[1699]) | (      i[1699]);
assign l_47[279]    = ( l_48 [133] & !i[1699]) | ( l_48 [144] &  i[1699]);
assign l_47[280]    = ( l_48 [145] & !i[1699]) | (      i[1699]);
assign l_47[281]    = ( l_48 [133] & !i[1699]) | ( l_48 [145] &  i[1699]);
assign l_47[282]    = ( l_48 [146] & !i[1699]) | (      i[1699]);
assign l_47[283]    = ( l_48 [133] & !i[1699]) | ( l_48 [146] &  i[1699]);
assign l_47[284]    = ( l_48 [147] & !i[1699]) | (      i[1699]);
assign l_47[285]    = ( l_48 [133] & !i[1699]) | ( l_48 [147] &  i[1699]);
assign l_47[286]    = ( l_48 [148] & !i[1699]) | (      i[1699]);
assign l_47[287]    = ( l_48 [133] & !i[1699]) | ( l_48 [148] &  i[1699]);
assign l_47[288]    = ( l_48 [149] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[289]    = ( l_48 [150] & !i[1699]) | ( l_48 [149] &  i[1699]);
assign l_47[290]    = ( l_48 [151] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[291]    = ( l_48 [150] & !i[1699]) | ( l_48 [151] &  i[1699]);
assign l_47[292]    = ( l_48 [152] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[293]    = ( l_48 [150] & !i[1699]) | ( l_48 [152] &  i[1699]);
assign l_47[294]    = ( l_48 [153] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[295]    = ( l_48 [150] & !i[1699]) | ( l_48 [153] &  i[1699]);
assign l_47[296]    = ( l_48 [154] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[297]    = ( l_48 [150] & !i[1699]) | ( l_48 [154] &  i[1699]);
assign l_47[298]    = ( l_48 [155] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[299]    = ( l_48 [150] & !i[1699]) | ( l_48 [155] &  i[1699]);
assign l_47[300]    = ( l_48 [156] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[301]    = ( l_48 [150] & !i[1699]) | ( l_48 [156] &  i[1699]);
assign l_47[302]    = ( l_48 [157] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[303]    = ( l_48 [150] & !i[1699]) | ( l_48 [157] &  i[1699]);
assign l_47[304]    = ( l_48 [158] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[305]    = ( l_48 [150] & !i[1699]) | ( l_48 [158] &  i[1699]);
assign l_47[306]    = ( l_48 [159] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[307]    = ( l_48 [150] & !i[1699]) | ( l_48 [159] &  i[1699]);
assign l_47[308]    = ( l_48 [160] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[309]    = ( l_48 [150] & !i[1699]) | ( l_48 [160] &  i[1699]);
assign l_47[310]    = ( l_48 [161] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[311]    = ( l_48 [150] & !i[1699]) | ( l_48 [161] &  i[1699]);
assign l_47[312]    = ( l_48 [162] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[313]    = ( l_48 [150] & !i[1699]) | ( l_48 [162] &  i[1699]);
assign l_47[314]    = ( l_48 [163] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[315]    = ( l_48 [150] & !i[1699]) | ( l_48 [163] &  i[1699]);
assign l_47[316]    = ( l_48 [164] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[317]    = ( l_48 [150] & !i[1699]) | ( l_48 [164] &  i[1699]);
assign l_47[318]    = ( l_48 [165] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[319]    = ( l_48 [150] & !i[1699]) | ( l_48 [165] &  i[1699]);
assign l_47[320]    = ( l_48 [166] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[321]    = ( l_48 [167] & !i[1699]) | ( l_48 [166] &  i[1699]);
assign l_47[322]    = ( l_48 [168] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[323]    = ( l_48 [167] & !i[1699]) | ( l_48 [168] &  i[1699]);
assign l_47[324]    = ( l_48 [169] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[325]    = ( l_48 [167] & !i[1699]) | ( l_48 [169] &  i[1699]);
assign l_47[326]    = ( l_48 [170] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[327]    = ( l_48 [167] & !i[1699]) | ( l_48 [170] &  i[1699]);
assign l_47[328]    = ( l_48 [171] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[329]    = ( l_48 [167] & !i[1699]) | ( l_48 [171] &  i[1699]);
assign l_47[330]    = ( l_48 [172] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[331]    = ( l_48 [167] & !i[1699]) | ( l_48 [172] &  i[1699]);
assign l_47[332]    = ( l_48 [173] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[333]    = ( l_48 [167] & !i[1699]) | ( l_48 [173] &  i[1699]);
assign l_47[334]    = ( l_48 [174] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[335]    = ( l_48 [167] & !i[1699]) | ( l_48 [174] &  i[1699]);
assign l_47[336]    = ( l_48 [175] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[337]    = ( l_48 [167] & !i[1699]) | ( l_48 [175] &  i[1699]);
assign l_47[338]    = ( l_48 [176] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[339]    = ( l_48 [167] & !i[1699]) | ( l_48 [176] &  i[1699]);
assign l_47[340]    = ( l_48 [177] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[341]    = ( l_48 [167] & !i[1699]) | ( l_48 [177] &  i[1699]);
assign l_47[342]    = ( l_48 [178] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[343]    = ( l_48 [167] & !i[1699]) | ( l_48 [178] &  i[1699]);
assign l_47[344]    = ( l_48 [179] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[345]    = ( l_48 [167] & !i[1699]) | ( l_48 [179] &  i[1699]);
assign l_47[346]    = ( l_48 [180] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[347]    = ( l_48 [167] & !i[1699]) | ( l_48 [180] &  i[1699]);
assign l_47[348]    = ( l_48 [181] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[349]    = ( l_48 [167] & !i[1699]) | ( l_48 [181] &  i[1699]);
assign l_47[350]    = ( l_48 [182] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[351]    = ( l_48 [167] & !i[1699]) | ( l_48 [182] &  i[1699]);
assign l_47[352]    = ( l_48 [183] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[353]    = ( l_48 [1] & !i[1699]) | ( l_48 [183] &  i[1699]);
assign l_47[354]    = ( l_48 [184] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[355]    = ( l_48 [1] & !i[1699]) | ( l_48 [184] &  i[1699]);
assign l_47[356]    = ( l_48 [185] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[357]    = ( l_48 [1] & !i[1699]) | ( l_48 [185] &  i[1699]);
assign l_47[358]    = ( l_48 [186] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[359]    = ( l_48 [1] & !i[1699]) | ( l_48 [186] &  i[1699]);
assign l_47[360]    = ( l_48 [187] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[361]    = ( l_48 [1] & !i[1699]) | ( l_48 [187] &  i[1699]);
assign l_47[362]    = ( l_48 [188] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[363]    = ( l_48 [1] & !i[1699]) | ( l_48 [188] &  i[1699]);
assign l_47[364]    = ( l_48 [189] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[365]    = ( l_48 [1] & !i[1699]) | ( l_48 [189] &  i[1699]);
assign l_47[366]    = ( l_48 [190] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[367]    = ( l_48 [1] & !i[1699]) | ( l_48 [190] &  i[1699]);
assign l_47[368]    = ( l_48 [191] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[369]    = ( l_48 [1] & !i[1699]) | ( l_48 [191] &  i[1699]);
assign l_47[370]    = ( l_48 [192] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[371]    = ( l_48 [1] & !i[1699]) | ( l_48 [192] &  i[1699]);
assign l_47[372]    = ( l_48 [193] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[373]    = ( l_48 [1] & !i[1699]) | ( l_48 [193] &  i[1699]);
assign l_47[374]    = ( l_48 [194] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[375]    = ( l_48 [1] & !i[1699]) | ( l_48 [194] &  i[1699]);
assign l_47[376]    = ( l_48 [195] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[377]    = ( l_48 [1] & !i[1699]) | ( l_48 [195] &  i[1699]);
assign l_47[378]    = ( l_48 [196] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[379]    = ( l_48 [1] & !i[1699]) | ( l_48 [196] &  i[1699]);
assign l_47[380]    = ( l_48 [197] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[381]    = ( l_48 [1] & !i[1699]) | ( l_48 [197] &  i[1699]);
assign l_47[382]    = ( l_48 [198] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[383]    = ( l_48 [1] & !i[1699]) | ( l_48 [198] &  i[1699]);
assign l_47[384]    = ( l_48 [199] & !i[1699]) | (      i[1699]);
assign l_47[385]    = ( l_48 [133] & !i[1699]) | ( l_48 [199] &  i[1699]);
assign l_47[386]    = ( l_48 [200] & !i[1699]) | (      i[1699]);
assign l_47[387]    = ( l_48 [133] & !i[1699]) | ( l_48 [200] &  i[1699]);
assign l_47[388]    = ( l_48 [201] & !i[1699]) | (      i[1699]);
assign l_47[389]    = ( l_48 [133] & !i[1699]) | ( l_48 [201] &  i[1699]);
assign l_47[390]    = ( l_48 [202] & !i[1699]) | (      i[1699]);
assign l_47[391]    = ( l_48 [133] & !i[1699]) | ( l_48 [202] &  i[1699]);
assign l_47[392]    = ( l_48 [203] & !i[1699]) | (      i[1699]);
assign l_47[393]    = ( l_48 [133] & !i[1699]) | ( l_48 [203] &  i[1699]);
assign l_47[394]    = ( l_48 [204] & !i[1699]) | (      i[1699]);
assign l_47[395]    = ( l_48 [133] & !i[1699]) | ( l_48 [204] &  i[1699]);
assign l_47[396]    = ( l_48 [205] & !i[1699]) | (      i[1699]);
assign l_47[397]    = ( l_48 [133] & !i[1699]) | ( l_48 [205] &  i[1699]);
assign l_47[398]    = ( l_48 [206] & !i[1699]) | (      i[1699]);
assign l_47[399]    = ( l_48 [133] & !i[1699]) | ( l_48 [206] &  i[1699]);
assign l_47[400]    = ( l_48 [207] & !i[1699]) | (      i[1699]);
assign l_47[401]    = ( l_48 [133] & !i[1699]) | ( l_48 [207] &  i[1699]);
assign l_47[402]    = ( l_48 [208] & !i[1699]) | (      i[1699]);
assign l_47[403]    = ( l_48 [133] & !i[1699]) | ( l_48 [208] &  i[1699]);
assign l_47[404]    = ( l_48 [209] & !i[1699]) | (      i[1699]);
assign l_47[405]    = ( l_48 [133] & !i[1699]) | ( l_48 [209] &  i[1699]);
assign l_47[406]    = ( l_48 [210] & !i[1699]) | (      i[1699]);
assign l_47[407]    = ( l_48 [133] & !i[1699]) | ( l_48 [210] &  i[1699]);
assign l_47[408]    = ( l_48 [211] & !i[1699]) | (      i[1699]);
assign l_47[409]    = ( l_48 [133] & !i[1699]) | ( l_48 [211] &  i[1699]);
assign l_47[410]    = ( l_48 [212] & !i[1699]) | (      i[1699]);
assign l_47[411]    = ( l_48 [133] & !i[1699]) | ( l_48 [212] &  i[1699]);
assign l_47[412]    = ( l_48 [213] & !i[1699]) | (      i[1699]);
assign l_47[413]    = ( l_48 [133] & !i[1699]) | ( l_48 [213] &  i[1699]);
assign l_47[414]    = ( l_48 [214] & !i[1699]) | (      i[1699]);
assign l_47[415]    = ( l_48 [133] & !i[1699]) | ( l_48 [214] &  i[1699]);
assign l_47[416]    = ( l_48 [215] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[417]    = ( l_48 [150] & !i[1699]) | ( l_48 [215] &  i[1699]);
assign l_47[418]    = ( l_48 [216] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[419]    = ( l_48 [150] & !i[1699]) | ( l_48 [216] &  i[1699]);
assign l_47[420]    = ( l_48 [217] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[421]    = ( l_48 [150] & !i[1699]) | ( l_48 [217] &  i[1699]);
assign l_47[422]    = ( l_48 [218] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[423]    = ( l_48 [150] & !i[1699]) | ( l_48 [218] &  i[1699]);
assign l_47[424]    = ( l_48 [219] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[425]    = ( l_48 [150] & !i[1699]) | ( l_48 [219] &  i[1699]);
assign l_47[426]    = ( l_48 [220] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[427]    = ( l_48 [150] & !i[1699]) | ( l_48 [220] &  i[1699]);
assign l_47[428]    = ( l_48 [221] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[429]    = ( l_48 [150] & !i[1699]) | ( l_48 [221] &  i[1699]);
assign l_47[430]    = ( l_48 [222] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[431]    = ( l_48 [150] & !i[1699]) | ( l_48 [222] &  i[1699]);
assign l_47[432]    = ( l_48 [223] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[433]    = ( l_48 [150] & !i[1699]) | ( l_48 [223] &  i[1699]);
assign l_47[434]    = ( l_48 [224] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[435]    = ( l_48 [150] & !i[1699]) | ( l_48 [224] &  i[1699]);
assign l_47[436]    = ( l_48 [225] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[437]    = ( l_48 [150] & !i[1699]) | ( l_48 [225] &  i[1699]);
assign l_47[438]    = ( l_48 [226] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[439]    = ( l_48 [150] & !i[1699]) | ( l_48 [226] &  i[1699]);
assign l_47[440]    = ( l_48 [227] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[441]    = ( l_48 [150] & !i[1699]) | ( l_48 [227] &  i[1699]);
assign l_47[442]    = ( l_48 [228] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[443]    = ( l_48 [150] & !i[1699]) | ( l_48 [228] &  i[1699]);
assign l_47[444]    = ( l_48 [229] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[445]    = ( l_48 [150] & !i[1699]) | ( l_48 [229] &  i[1699]);
assign l_47[446]    = ( l_48 [230] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[447]    = ( l_48 [150] & !i[1699]) | ( l_48 [230] &  i[1699]);
assign l_47[448]    = ( l_48 [231] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[449]    = ( l_48 [167] & !i[1699]) | ( l_48 [231] &  i[1699]);
assign l_47[450]    = ( l_48 [232] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[451]    = ( l_48 [167] & !i[1699]) | ( l_48 [232] &  i[1699]);
assign l_47[452]    = ( l_48 [233] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[453]    = ( l_48 [167] & !i[1699]) | ( l_48 [233] &  i[1699]);
assign l_47[454]    = ( l_48 [234] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[455]    = ( l_48 [167] & !i[1699]) | ( l_48 [234] &  i[1699]);
assign l_47[456]    = ( l_48 [235] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[457]    = ( l_48 [167] & !i[1699]) | ( l_48 [235] &  i[1699]);
assign l_47[458]    = ( l_48 [236] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[459]    = ( l_48 [167] & !i[1699]) | ( l_48 [236] &  i[1699]);
assign l_47[460]    = ( l_48 [237] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[461]    = ( l_48 [167] & !i[1699]) | ( l_48 [237] &  i[1699]);
assign l_47[462]    = ( l_48 [238] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[463]    = ( l_48 [167] & !i[1699]) | ( l_48 [238] &  i[1699]);
assign l_47[464]    = ( l_48 [239] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[465]    = ( l_48 [167] & !i[1699]) | ( l_48 [239] &  i[1699]);
assign l_47[466]    = ( l_48 [240] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[467]    = ( l_48 [167] & !i[1699]) | ( l_48 [240] &  i[1699]);
assign l_47[468]    = ( l_48 [241] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[469]    = ( l_48 [167] & !i[1699]) | ( l_48 [241] &  i[1699]);
assign l_47[470]    = ( l_48 [242] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[471]    = ( l_48 [167] & !i[1699]) | ( l_48 [242] &  i[1699]);
assign l_47[472]    = ( l_48 [243] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[473]    = ( l_48 [167] & !i[1699]) | ( l_48 [243] &  i[1699]);
assign l_47[474]    = ( l_48 [244] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[475]    = ( l_48 [167] & !i[1699]) | ( l_48 [244] &  i[1699]);
assign l_47[476]    = ( l_48 [245] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[477]    = ( l_48 [167] & !i[1699]) | ( l_48 [245] &  i[1699]);
assign l_47[478]    = ( l_48 [246] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[479]    = ( l_48 [167] & !i[1699]) | ( l_48 [246] &  i[1699]);
assign l_47[480]    = ( l_48 [247] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[481]    = ( l_48 [1] & !i[1699]) | ( l_48 [247] &  i[1699]);
assign l_47[482]    = ( l_48 [248] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[483]    = ( l_48 [1] & !i[1699]) | ( l_48 [248] &  i[1699]);
assign l_47[484]    = ( l_48 [249] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[485]    = ( l_48 [1] & !i[1699]) | ( l_48 [249] &  i[1699]);
assign l_47[486]    = ( l_48 [250] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[487]    = ( l_48 [1] & !i[1699]) | ( l_48 [250] &  i[1699]);
assign l_47[488]    = ( l_48 [251] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[489]    = ( l_48 [1] & !i[1699]) | ( l_48 [251] &  i[1699]);
assign l_47[490]    = ( l_48 [252] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[491]    = ( l_48 [1] & !i[1699]) | ( l_48 [252] &  i[1699]);
assign l_47[492]    = ( l_48 [253] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[493]    = ( l_48 [1] & !i[1699]) | ( l_48 [253] &  i[1699]);
assign l_47[494]    = ( l_48 [254] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[495]    = ( l_48 [1] & !i[1699]) | ( l_48 [254] &  i[1699]);
assign l_47[496]    = ( l_48 [255] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[497]    = ( l_48 [1] & !i[1699]) | ( l_48 [255] &  i[1699]);
assign l_47[498]    = ( l_48 [256] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[499]    = ( l_48 [1] & !i[1699]) | ( l_48 [256] &  i[1699]);
assign l_47[500]    = ( l_48 [257] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[501]    = ( l_48 [1] & !i[1699]) | ( l_48 [257] &  i[1699]);
assign l_47[502]    = ( l_48 [258] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[503]    = ( l_48 [1] & !i[1699]) | ( l_48 [258] &  i[1699]);
assign l_47[504]    = ( l_48 [259] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[505]    = ( l_48 [1] & !i[1699]) | ( l_48 [259] &  i[1699]);
assign l_47[506]    = ( l_48 [260] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[507]    = ( l_48 [1] & !i[1699]) | ( l_48 [260] &  i[1699]);
assign l_47[508]    = ( l_48 [261] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[509]    = ( l_48 [1] & !i[1699]) | ( l_48 [261] &  i[1699]);
assign l_47[510]    = ( l_48 [262] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[511]    = ( l_48 [1] & !i[1699]) | ( l_48 [262] &  i[1699]);
assign l_47[512]    = ( l_48 [263] & !i[1699]) | ( l_48 [1] &  i[1699]);
assign l_47[513]    = ( l_48 [2] & !i[1699]) | ( l_48 [263] &  i[1699]);
assign l_47[514]    = ( l_48 [264] & !i[1699]) | ( l_48 [2] &  i[1699]);
assign l_47[515]    = ( l_48 [19] & !i[1699]) | ( l_48 [264] &  i[1699]);
assign l_47[516]    = ( l_48 [265] & !i[1699]) | ( l_48 [19] &  i[1699]);
assign l_47[517]    = ( l_48 [36] & !i[1699]) | ( l_48 [265] &  i[1699]);
assign l_47[518]    = ( l_48 [266] & !i[1699]) | ( l_48 [36] &  i[1699]);
assign l_47[519]    = ( l_48 [266] &  i[1699]);
assign l_47[520]    = ( l_48 [267] & !i[1699]) | (      i[1699]);
assign l_47[521]    = ( l_48 [133] & !i[1699]) | ( l_48 [267] &  i[1699]);
assign l_47[522]    = ( l_48 [268] & !i[1699]) | ( l_48 [133] &  i[1699]);
assign l_47[523]    = ( l_48 [150] & !i[1699]) | ( l_48 [268] &  i[1699]);
assign l_47[524]    = ( l_48 [269] & !i[1699]) | ( l_48 [150] &  i[1699]);
assign l_47[525]    = ( l_48 [167] & !i[1699]) | ( l_48 [269] &  i[1699]);
assign l_47[526]    = ( l_48 [270] & !i[1699]) | ( l_48 [167] &  i[1699]);
assign l_47[527]    = ( l_48 [1] & !i[1699]) | ( l_48 [270] &  i[1699]);
assign l_47[528]    = ( l_48 [271] & !i[1699]) | (      i[1699]);
assign l_47[529]    = ( l_48 [272] & !i[1699]) | ( l_48 [271] &  i[1699]);
assign l_47[530]    = ( l_48 [273] & !i[1699]) | (      i[1699]);
assign l_47[531]    = ( l_48 [272] & !i[1699]) | ( l_48 [273] &  i[1699]);
assign l_47[532]    = ( l_48 [274] & !i[1699]) | (      i[1699]);
assign l_47[533]    = ( l_48 [272] & !i[1699]) | ( l_48 [274] &  i[1699]);
assign l_47[534]    = ( l_48 [275] & !i[1699]) | (      i[1699]);
assign l_47[535]    = ( l_48 [272] & !i[1699]) | ( l_48 [275] &  i[1699]);
assign l_47[536]    = ( l_48 [276] & !i[1699]) | (      i[1699]);
assign l_47[537]    = ( l_48 [272] & !i[1699]) | ( l_48 [276] &  i[1699]);
assign l_47[538]    = ( l_48 [277] & !i[1699]) | (      i[1699]);
assign l_47[539]    = ( l_48 [272] & !i[1699]) | ( l_48 [277] &  i[1699]);
assign l_47[540]    = ( l_48 [278] & !i[1699]) | (      i[1699]);
assign l_47[541]    = ( l_48 [272] & !i[1699]) | ( l_48 [278] &  i[1699]);
assign l_47[542]    = ( l_48 [279] & !i[1699]) | (      i[1699]);
assign l_47[543]    = ( l_48 [272] & !i[1699]) | ( l_48 [279] &  i[1699]);
assign l_47[544]    = ( l_48 [280] & !i[1699]) | (      i[1699]);
assign l_47[545]    = ( l_48 [272] & !i[1699]) | ( l_48 [280] &  i[1699]);
assign l_47[546]    = ( l_48 [281] & !i[1699]) | (      i[1699]);
assign l_47[547]    = ( l_48 [272] & !i[1699]) | ( l_48 [281] &  i[1699]);
assign l_47[548]    = ( l_48 [282] & !i[1699]) | (      i[1699]);
assign l_47[549]    = ( l_48 [272] & !i[1699]) | ( l_48 [282] &  i[1699]);
assign l_47[550]    = ( l_48 [283] & !i[1699]) | (      i[1699]);
assign l_47[551]    = ( l_48 [272] & !i[1699]) | ( l_48 [283] &  i[1699]);
assign l_47[552]    = ( l_48 [284] & !i[1699]) | (      i[1699]);
assign l_47[553]    = ( l_48 [272] & !i[1699]) | ( l_48 [284] &  i[1699]);
assign l_47[554]    = ( l_48 [285] & !i[1699]) | (      i[1699]);
assign l_47[555]    = ( l_48 [272] & !i[1699]) | ( l_48 [285] &  i[1699]);
assign l_47[556]    = ( l_48 [286] & !i[1699]) | (      i[1699]);
assign l_47[557]    = ( l_48 [272] & !i[1699]) | ( l_48 [286] &  i[1699]);
assign l_47[558]    = ( l_48 [287] & !i[1699]) | (      i[1699]);
assign l_47[559]    = ( l_48 [272] & !i[1699]) | ( l_48 [287] &  i[1699]);
assign l_47[560]    = ( l_48 [288] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[561]    = ( l_48 [289] & !i[1699]) | ( l_48 [288] &  i[1699]);
assign l_47[562]    = ( l_48 [290] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[563]    = ( l_48 [289] & !i[1699]) | ( l_48 [290] &  i[1699]);
assign l_47[564]    = ( l_48 [291] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[565]    = ( l_48 [289] & !i[1699]) | ( l_48 [291] &  i[1699]);
assign l_47[566]    = ( l_48 [292] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[567]    = ( l_48 [289] & !i[1699]) | ( l_48 [292] &  i[1699]);
assign l_47[568]    = ( l_48 [293] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[569]    = ( l_48 [289] & !i[1699]) | ( l_48 [293] &  i[1699]);
assign l_47[570]    = ( l_48 [294] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[571]    = ( l_48 [289] & !i[1699]) | ( l_48 [294] &  i[1699]);
assign l_47[572]    = ( l_48 [295] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[573]    = ( l_48 [289] & !i[1699]) | ( l_48 [295] &  i[1699]);
assign l_47[574]    = ( l_48 [296] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[575]    = ( l_48 [289] & !i[1699]) | ( l_48 [296] &  i[1699]);
assign l_47[576]    = ( l_48 [297] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[577]    = ( l_48 [289] & !i[1699]) | ( l_48 [297] &  i[1699]);
assign l_47[578]    = ( l_48 [298] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[579]    = ( l_48 [289] & !i[1699]) | ( l_48 [298] &  i[1699]);
assign l_47[580]    = ( l_48 [299] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[581]    = ( l_48 [289] & !i[1699]) | ( l_48 [299] &  i[1699]);
assign l_47[582]    = ( l_48 [300] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[583]    = ( l_48 [289] & !i[1699]) | ( l_48 [300] &  i[1699]);
assign l_47[584]    = ( l_48 [301] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[585]    = ( l_48 [289] & !i[1699]) | ( l_48 [301] &  i[1699]);
assign l_47[586]    = ( l_48 [302] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[587]    = ( l_48 [289] & !i[1699]) | ( l_48 [302] &  i[1699]);
assign l_47[588]    = ( l_48 [303] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[589]    = ( l_48 [289] & !i[1699]) | ( l_48 [303] &  i[1699]);
assign l_47[590]    = ( l_48 [304] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[591]    = ( l_48 [289] & !i[1699]) | ( l_48 [304] &  i[1699]);
assign l_47[592]    = ( l_48 [305] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[593]    = ( l_48 [306] & !i[1699]) | ( l_48 [305] &  i[1699]);
assign l_47[594]    = ( l_48 [307] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[595]    = ( l_48 [306] & !i[1699]) | ( l_48 [307] &  i[1699]);
assign l_47[596]    = ( l_48 [308] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[597]    = ( l_48 [306] & !i[1699]) | ( l_48 [308] &  i[1699]);
assign l_47[598]    = ( l_48 [309] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[599]    = ( l_48 [306] & !i[1699]) | ( l_48 [309] &  i[1699]);
assign l_47[600]    = ( l_48 [310] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[601]    = ( l_48 [306] & !i[1699]) | ( l_48 [310] &  i[1699]);
assign l_47[602]    = ( l_48 [311] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[603]    = ( l_48 [306] & !i[1699]) | ( l_48 [311] &  i[1699]);
assign l_47[604]    = ( l_48 [312] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[605]    = ( l_48 [306] & !i[1699]) | ( l_48 [312] &  i[1699]);
assign l_47[606]    = ( l_48 [313] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[607]    = ( l_48 [306] & !i[1699]) | ( l_48 [313] &  i[1699]);
assign l_47[608]    = ( l_48 [314] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[609]    = ( l_48 [306] & !i[1699]) | ( l_48 [314] &  i[1699]);
assign l_47[610]    = ( l_48 [315] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[611]    = ( l_48 [306] & !i[1699]) | ( l_48 [315] &  i[1699]);
assign l_47[612]    = ( l_48 [316] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[613]    = ( l_48 [306] & !i[1699]) | ( l_48 [316] &  i[1699]);
assign l_47[614]    = ( l_48 [317] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[615]    = ( l_48 [306] & !i[1699]) | ( l_48 [317] &  i[1699]);
assign l_47[616]    = ( l_48 [318] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[617]    = ( l_48 [306] & !i[1699]) | ( l_48 [318] &  i[1699]);
assign l_47[618]    = ( l_48 [319] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[619]    = ( l_48 [306] & !i[1699]) | ( l_48 [319] &  i[1699]);
assign l_47[620]    = ( l_48 [320] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[621]    = ( l_48 [306] & !i[1699]) | ( l_48 [320] &  i[1699]);
assign l_47[622]    = ( l_48 [321] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[623]    = ( l_48 [306] & !i[1699]) | ( l_48 [321] &  i[1699]);
assign l_47[624]    = ( l_48 [322] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[625]    = (!l_48 [1] & !i[1699]) | ( l_48 [322] &  i[1699]);
assign l_47[626]    = ( l_48 [323] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[627]    = (!l_48 [1] & !i[1699]) | ( l_48 [323] &  i[1699]);
assign l_47[628]    = ( l_48 [324] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[629]    = (!l_48 [1] & !i[1699]) | ( l_48 [324] &  i[1699]);
assign l_47[630]    = ( l_48 [325] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[631]    = (!l_48 [1] & !i[1699]) | ( l_48 [325] &  i[1699]);
assign l_47[632]    = ( l_48 [326] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[633]    = (!l_48 [1] & !i[1699]) | ( l_48 [326] &  i[1699]);
assign l_47[634]    = ( l_48 [327] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[635]    = (!l_48 [1] & !i[1699]) | ( l_48 [327] &  i[1699]);
assign l_47[636]    = ( l_48 [328] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[637]    = (!l_48 [1] & !i[1699]) | ( l_48 [328] &  i[1699]);
assign l_47[638]    = ( l_48 [329] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[639]    = (!l_48 [1] & !i[1699]) | ( l_48 [329] &  i[1699]);
assign l_47[640]    = ( l_48 [330] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[641]    = (!l_48 [1] & !i[1699]) | ( l_48 [330] &  i[1699]);
assign l_47[642]    = ( l_48 [331] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[643]    = (!l_48 [1] & !i[1699]) | ( l_48 [331] &  i[1699]);
assign l_47[644]    = ( l_48 [332] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[645]    = (!l_48 [1] & !i[1699]) | ( l_48 [332] &  i[1699]);
assign l_47[646]    = ( l_48 [333] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[647]    = (!l_48 [1] & !i[1699]) | ( l_48 [333] &  i[1699]);
assign l_47[648]    = ( l_48 [334] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[649]    = (!l_48 [1] & !i[1699]) | ( l_48 [334] &  i[1699]);
assign l_47[650]    = ( l_48 [335] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[651]    = (!l_48 [1] & !i[1699]) | ( l_48 [335] &  i[1699]);
assign l_47[652]    = ( l_48 [336] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[653]    = (!l_48 [1] & !i[1699]) | ( l_48 [336] &  i[1699]);
assign l_47[654]    = ( l_48 [337] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[655]    = (!l_48 [1] & !i[1699]) | ( l_48 [337] &  i[1699]);
assign l_47[656]    = (!l_48 [1] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[657]    = ( l_48 [339] & !i[1699]) | (      i[1699]);
assign l_47[658]    = ( l_48 [272] & !i[1699]) | ( l_48 [339] &  i[1699]);
assign l_47[659]    = ( l_48 [340] & !i[1699]) | (      i[1699]);
assign l_47[660]    = ( l_48 [272] & !i[1699]) | ( l_48 [340] &  i[1699]);
assign l_47[661]    = ( l_48 [341] & !i[1699]) | (      i[1699]);
assign l_47[662]    = ( l_48 [272] & !i[1699]) | ( l_48 [341] &  i[1699]);
assign l_47[663]    = ( l_48 [342] & !i[1699]) | (      i[1699]);
assign l_47[664]    = ( l_48 [272] & !i[1699]) | ( l_48 [342] &  i[1699]);
assign l_47[665]    = ( l_48 [343] & !i[1699]) | (      i[1699]);
assign l_47[666]    = ( l_48 [272] & !i[1699]) | ( l_48 [343] &  i[1699]);
assign l_47[667]    = ( l_48 [344] & !i[1699]) | (      i[1699]);
assign l_47[668]    = ( l_48 [272] & !i[1699]) | ( l_48 [344] &  i[1699]);
assign l_47[669]    = ( l_48 [345] & !i[1699]) | (      i[1699]);
assign l_47[670]    = ( l_48 [272] & !i[1699]) | ( l_48 [345] &  i[1699]);
assign l_47[671]    = ( l_48 [346] & !i[1699]) | (      i[1699]);
assign l_47[672]    = ( l_48 [272] & !i[1699]) | ( l_48 [346] &  i[1699]);
assign l_47[673]    = ( l_48 [347] & !i[1699]) | (      i[1699]);
assign l_47[674]    = ( l_48 [272] & !i[1699]) | ( l_48 [347] &  i[1699]);
assign l_47[675]    = ( l_48 [348] & !i[1699]) | (      i[1699]);
assign l_47[676]    = ( l_48 [272] & !i[1699]) | ( l_48 [348] &  i[1699]);
assign l_47[677]    = ( l_48 [349] & !i[1699]) | (      i[1699]);
assign l_47[678]    = ( l_48 [272] & !i[1699]) | ( l_48 [349] &  i[1699]);
assign l_47[679]    = ( l_48 [350] & !i[1699]) | (      i[1699]);
assign l_47[680]    = ( l_48 [272] & !i[1699]) | ( l_48 [350] &  i[1699]);
assign l_47[681]    = ( l_48 [351] & !i[1699]) | (      i[1699]);
assign l_47[682]    = ( l_48 [272] & !i[1699]) | ( l_48 [351] &  i[1699]);
assign l_47[683]    = ( l_48 [352] & !i[1699]) | (      i[1699]);
assign l_47[684]    = ( l_48 [272] & !i[1699]) | ( l_48 [352] &  i[1699]);
assign l_47[685]    = ( l_48 [353] & !i[1699]) | (      i[1699]);
assign l_47[686]    = ( l_48 [272] & !i[1699]) | ( l_48 [353] &  i[1699]);
assign l_47[687]    = ( l_48 [354] & !i[1699]) | (      i[1699]);
assign l_47[688]    = ( l_48 [272] & !i[1699]) | ( l_48 [354] &  i[1699]);
assign l_47[689]    = ( l_48 [355] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[690]    = ( l_48 [289] & !i[1699]) | ( l_48 [355] &  i[1699]);
assign l_47[691]    = ( l_48 [356] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[692]    = ( l_48 [289] & !i[1699]) | ( l_48 [356] &  i[1699]);
assign l_47[693]    = ( l_48 [357] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[694]    = ( l_48 [289] & !i[1699]) | ( l_48 [357] &  i[1699]);
assign l_47[695]    = ( l_48 [358] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[696]    = ( l_48 [289] & !i[1699]) | ( l_48 [358] &  i[1699]);
assign l_47[697]    = ( l_48 [359] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[698]    = ( l_48 [289] & !i[1699]) | ( l_48 [359] &  i[1699]);
assign l_47[699]    = ( l_48 [360] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[700]    = ( l_48 [289] & !i[1699]) | ( l_48 [360] &  i[1699]);
assign l_47[701]    = ( l_48 [361] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[702]    = ( l_48 [289] & !i[1699]) | ( l_48 [361] &  i[1699]);
assign l_47[703]    = ( l_48 [362] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[704]    = ( l_48 [289] & !i[1699]) | ( l_48 [362] &  i[1699]);
assign l_47[705]    = ( l_48 [363] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[706]    = ( l_48 [289] & !i[1699]) | ( l_48 [363] &  i[1699]);
assign l_47[707]    = ( l_48 [364] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[708]    = ( l_48 [289] & !i[1699]) | ( l_48 [364] &  i[1699]);
assign l_47[709]    = ( l_48 [365] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[710]    = ( l_48 [289] & !i[1699]) | ( l_48 [365] &  i[1699]);
assign l_47[711]    = ( l_48 [366] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[712]    = ( l_48 [289] & !i[1699]) | ( l_48 [366] &  i[1699]);
assign l_47[713]    = ( l_48 [367] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[714]    = ( l_48 [289] & !i[1699]) | ( l_48 [367] &  i[1699]);
assign l_47[715]    = ( l_48 [368] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[716]    = ( l_48 [289] & !i[1699]) | ( l_48 [368] &  i[1699]);
assign l_47[717]    = ( l_48 [369] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[718]    = ( l_48 [289] & !i[1699]) | ( l_48 [369] &  i[1699]);
assign l_47[719]    = ( l_48 [370] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[720]    = ( l_48 [289] & !i[1699]) | ( l_48 [370] &  i[1699]);
assign l_47[721]    = ( l_48 [371] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[722]    = ( l_48 [306] & !i[1699]) | ( l_48 [371] &  i[1699]);
assign l_47[723]    = ( l_48 [372] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[724]    = ( l_48 [306] & !i[1699]) | ( l_48 [372] &  i[1699]);
assign l_47[725]    = ( l_48 [373] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[726]    = ( l_48 [306] & !i[1699]) | ( l_48 [373] &  i[1699]);
assign l_47[727]    = ( l_48 [374] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[728]    = ( l_48 [306] & !i[1699]) | ( l_48 [374] &  i[1699]);
assign l_47[729]    = ( l_48 [375] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[730]    = ( l_48 [306] & !i[1699]) | ( l_48 [375] &  i[1699]);
assign l_47[731]    = ( l_48 [376] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[732]    = ( l_48 [306] & !i[1699]) | ( l_48 [376] &  i[1699]);
assign l_47[733]    = ( l_48 [377] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[734]    = ( l_48 [306] & !i[1699]) | ( l_48 [377] &  i[1699]);
assign l_47[735]    = ( l_48 [378] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[736]    = ( l_48 [306] & !i[1699]) | ( l_48 [378] &  i[1699]);
assign l_47[737]    = ( l_48 [379] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[738]    = ( l_48 [306] & !i[1699]) | ( l_48 [379] &  i[1699]);
assign l_47[739]    = ( l_48 [380] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[740]    = ( l_48 [306] & !i[1699]) | ( l_48 [380] &  i[1699]);
assign l_47[741]    = ( l_48 [381] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[742]    = ( l_48 [306] & !i[1699]) | ( l_48 [381] &  i[1699]);
assign l_47[743]    = ( l_48 [382] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[744]    = ( l_48 [306] & !i[1699]) | ( l_48 [382] &  i[1699]);
assign l_47[745]    = ( l_48 [383] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[746]    = ( l_48 [306] & !i[1699]) | ( l_48 [383] &  i[1699]);
assign l_47[747]    = ( l_48 [384] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[748]    = ( l_48 [306] & !i[1699]) | ( l_48 [384] &  i[1699]);
assign l_47[749]    = ( l_48 [385] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[750]    = ( l_48 [306] & !i[1699]) | ( l_48 [385] &  i[1699]);
assign l_47[751]    = ( l_48 [386] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[752]    = ( l_48 [306] & !i[1699]) | ( l_48 [386] &  i[1699]);
assign l_47[753]    = ( l_48 [387] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[754]    = ( l_48 [338] & !i[1699]) | ( l_48 [387] &  i[1699]);
assign l_47[755]    = ( l_48 [388] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[756]    = ( l_48 [338] & !i[1699]) | ( l_48 [388] &  i[1699]);
assign l_47[757]    = ( l_48 [389] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[758]    = ( l_48 [338] & !i[1699]) | ( l_48 [389] &  i[1699]);
assign l_47[759]    = ( l_48 [390] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[760]    = ( l_48 [338] & !i[1699]) | ( l_48 [390] &  i[1699]);
assign l_47[761]    = ( l_48 [391] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[762]    = ( l_48 [338] & !i[1699]) | ( l_48 [391] &  i[1699]);
assign l_47[763]    = ( l_48 [392] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[764]    = ( l_48 [338] & !i[1699]) | ( l_48 [392] &  i[1699]);
assign l_47[765]    = ( l_48 [393] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[766]    = ( l_48 [338] & !i[1699]) | ( l_48 [393] &  i[1699]);
assign l_47[767]    = ( l_48 [394] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[768]    = ( l_48 [338] & !i[1699]) | ( l_48 [394] &  i[1699]);
assign l_47[769]    = ( l_48 [395] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[770]    = ( l_48 [338] & !i[1699]) | ( l_48 [395] &  i[1699]);
assign l_47[771]    = ( l_48 [396] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[772]    = ( l_48 [338] & !i[1699]) | ( l_48 [396] &  i[1699]);
assign l_47[773]    = ( l_48 [397] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[774]    = ( l_48 [338] & !i[1699]) | ( l_48 [397] &  i[1699]);
assign l_47[775]    = ( l_48 [398] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[776]    = ( l_48 [338] & !i[1699]) | ( l_48 [398] &  i[1699]);
assign l_47[777]    = ( l_48 [399] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[778]    = ( l_48 [338] & !i[1699]) | ( l_48 [399] &  i[1699]);
assign l_47[779]    = ( l_48 [400] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[780]    = ( l_48 [338] & !i[1699]) | ( l_48 [400] &  i[1699]);
assign l_47[781]    = ( l_48 [401] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[782]    = ( l_48 [338] & !i[1699]) | ( l_48 [401] &  i[1699]);
assign l_47[783]    = ( l_48 [402] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[784]    = ( l_48 [338] & !i[1699]) | ( l_48 [402] &  i[1699]);
assign l_47[785]    = ( l_48 [403] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[786]    = ( l_48 [404] & !i[1699]) | ( l_48 [403] &  i[1699]);
assign l_47[787]    = ( l_48 [405] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[788]    = ( l_48 [404] & !i[1699]) | ( l_48 [405] &  i[1699]);
assign l_47[789]    = ( l_48 [406] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[790]    = ( l_48 [404] & !i[1699]) | ( l_48 [406] &  i[1699]);
assign l_47[791]    = ( l_48 [407] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[792]    = ( l_48 [404] & !i[1699]) | ( l_48 [407] &  i[1699]);
assign l_47[793]    = ( l_48 [408] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[794]    = ( l_48 [404] & !i[1699]) | ( l_48 [408] &  i[1699]);
assign l_47[795]    = ( l_48 [409] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[796]    = ( l_48 [404] & !i[1699]) | ( l_48 [409] &  i[1699]);
assign l_47[797]    = ( l_48 [410] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[798]    = ( l_48 [404] & !i[1699]) | ( l_48 [410] &  i[1699]);
assign l_47[799]    = ( l_48 [411] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[800]    = ( l_48 [404] & !i[1699]) | ( l_48 [411] &  i[1699]);
assign l_47[801]    = ( l_48 [412] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[802]    = ( l_48 [404] & !i[1699]) | ( l_48 [412] &  i[1699]);
assign l_47[803]    = ( l_48 [413] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[804]    = ( l_48 [404] & !i[1699]) | ( l_48 [413] &  i[1699]);
assign l_47[805]    = ( l_48 [414] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[806]    = ( l_48 [404] & !i[1699]) | ( l_48 [414] &  i[1699]);
assign l_47[807]    = ( l_48 [415] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[808]    = ( l_48 [404] & !i[1699]) | ( l_48 [415] &  i[1699]);
assign l_47[809]    = ( l_48 [416] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[810]    = ( l_48 [404] & !i[1699]) | ( l_48 [416] &  i[1699]);
assign l_47[811]    = ( l_48 [417] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[812]    = ( l_48 [404] & !i[1699]) | ( l_48 [417] &  i[1699]);
assign l_47[813]    = ( l_48 [418] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[814]    = ( l_48 [404] & !i[1699]) | ( l_48 [418] &  i[1699]);
assign l_47[815]    = ( l_48 [419] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[816]    = ( l_48 [404] & !i[1699]) | ( l_48 [419] &  i[1699]);
assign l_47[817]    = ( l_48 [420] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[818]    = ( l_48 [421] & !i[1699]) | ( l_48 [420] &  i[1699]);
assign l_47[819]    = ( l_48 [422] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[820]    = ( l_48 [421] & !i[1699]) | ( l_48 [422] &  i[1699]);
assign l_47[821]    = ( l_48 [423] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[822]    = ( l_48 [421] & !i[1699]) | ( l_48 [423] &  i[1699]);
assign l_47[823]    = ( l_48 [424] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[824]    = ( l_48 [421] & !i[1699]) | ( l_48 [424] &  i[1699]);
assign l_47[825]    = ( l_48 [425] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[826]    = ( l_48 [421] & !i[1699]) | ( l_48 [425] &  i[1699]);
assign l_47[827]    = ( l_48 [426] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[828]    = ( l_48 [421] & !i[1699]) | ( l_48 [426] &  i[1699]);
assign l_47[829]    = ( l_48 [427] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[830]    = ( l_48 [421] & !i[1699]) | ( l_48 [427] &  i[1699]);
assign l_47[831]    = ( l_48 [428] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[832]    = ( l_48 [421] & !i[1699]) | ( l_48 [428] &  i[1699]);
assign l_47[833]    = ( l_48 [429] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[834]    = ( l_48 [421] & !i[1699]) | ( l_48 [429] &  i[1699]);
assign l_47[835]    = ( l_48 [430] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[836]    = ( l_48 [421] & !i[1699]) | ( l_48 [430] &  i[1699]);
assign l_47[837]    = ( l_48 [431] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[838]    = ( l_48 [421] & !i[1699]) | ( l_48 [431] &  i[1699]);
assign l_47[839]    = ( l_48 [432] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[840]    = ( l_48 [421] & !i[1699]) | ( l_48 [432] &  i[1699]);
assign l_47[841]    = ( l_48 [433] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[842]    = ( l_48 [421] & !i[1699]) | ( l_48 [433] &  i[1699]);
assign l_47[843]    = ( l_48 [434] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[844]    = ( l_48 [421] & !i[1699]) | ( l_48 [434] &  i[1699]);
assign l_47[845]    = ( l_48 [435] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[846]    = ( l_48 [421] & !i[1699]) | ( l_48 [435] &  i[1699]);
assign l_47[847]    = ( l_48 [436] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[848]    = ( l_48 [421] & !i[1699]) | ( l_48 [436] &  i[1699]);
assign l_47[849]    = ( l_48 [437] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[850]    = ( l_48 [438] & !i[1699]) | ( l_48 [437] &  i[1699]);
assign l_47[851]    = ( l_48 [439] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[852]    = ( l_48 [438] & !i[1699]) | ( l_48 [439] &  i[1699]);
assign l_47[853]    = ( l_48 [440] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[854]    = ( l_48 [438] & !i[1699]) | ( l_48 [440] &  i[1699]);
assign l_47[855]    = ( l_48 [441] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[856]    = ( l_48 [438] & !i[1699]) | ( l_48 [441] &  i[1699]);
assign l_47[857]    = ( l_48 [442] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[858]    = ( l_48 [438] & !i[1699]) | ( l_48 [442] &  i[1699]);
assign l_47[859]    = ( l_48 [443] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[860]    = ( l_48 [438] & !i[1699]) | ( l_48 [443] &  i[1699]);
assign l_47[861]    = ( l_48 [444] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[862]    = ( l_48 [438] & !i[1699]) | ( l_48 [444] &  i[1699]);
assign l_47[863]    = ( l_48 [445] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[864]    = ( l_48 [438] & !i[1699]) | ( l_48 [445] &  i[1699]);
assign l_47[865]    = ( l_48 [446] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[866]    = ( l_48 [438] & !i[1699]) | ( l_48 [446] &  i[1699]);
assign l_47[867]    = ( l_48 [447] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[868]    = ( l_48 [438] & !i[1699]) | ( l_48 [447] &  i[1699]);
assign l_47[869]    = ( l_48 [448] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[870]    = ( l_48 [438] & !i[1699]) | ( l_48 [448] &  i[1699]);
assign l_47[871]    = ( l_48 [449] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[872]    = ( l_48 [438] & !i[1699]) | ( l_48 [449] &  i[1699]);
assign l_47[873]    = ( l_48 [450] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[874]    = ( l_48 [438] & !i[1699]) | ( l_48 [450] &  i[1699]);
assign l_47[875]    = ( l_48 [451] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[876]    = ( l_48 [438] & !i[1699]) | ( l_48 [451] &  i[1699]);
assign l_47[877]    = ( l_48 [452] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[878]    = ( l_48 [438] & !i[1699]) | ( l_48 [452] &  i[1699]);
assign l_47[879]    = ( l_48 [453] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[880]    = ( l_48 [438] & !i[1699]) | ( l_48 [453] &  i[1699]);
assign l_47[881]    = ( l_48 [454] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[882]    = ( l_48 [454] &  i[1699]);
assign l_47[883]    = ( l_48 [455] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[884]    = ( l_48 [455] &  i[1699]);
assign l_47[885]    = ( l_48 [456] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[886]    = ( l_48 [456] &  i[1699]);
assign l_47[887]    = ( l_48 [457] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[888]    = ( l_48 [457] &  i[1699]);
assign l_47[889]    = ( l_48 [458] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[890]    = ( l_48 [458] &  i[1699]);
assign l_47[891]    = ( l_48 [459] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[892]    = ( l_48 [459] &  i[1699]);
assign l_47[893]    = ( l_48 [460] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[894]    = ( l_48 [460] &  i[1699]);
assign l_47[895]    = ( l_48 [461] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[896]    = ( l_48 [461] &  i[1699]);
assign l_47[897]    = ( l_48 [462] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[898]    = ( l_48 [462] &  i[1699]);
assign l_47[899]    = ( l_48 [463] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[900]    = ( l_48 [463] &  i[1699]);
assign l_47[901]    = ( l_48 [464] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[902]    = ( l_48 [464] &  i[1699]);
assign l_47[903]    = ( l_48 [465] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[904]    = ( l_48 [465] &  i[1699]);
assign l_47[905]    = ( l_48 [466] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[906]    = ( l_48 [466] &  i[1699]);
assign l_47[907]    = ( l_48 [467] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[908]    = ( l_48 [467] &  i[1699]);
assign l_47[909]    = ( l_48 [468] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[910]    = ( l_48 [468] &  i[1699]);
assign l_47[911]    = ( l_48 [469] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[912]    = ( l_48 [469] &  i[1699]);
assign l_47[913]    = ( l_48 [470] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[914]    = ( l_48 [404] & !i[1699]) | ( l_48 [470] &  i[1699]);
assign l_47[915]    = ( l_48 [471] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[916]    = ( l_48 [404] & !i[1699]) | ( l_48 [471] &  i[1699]);
assign l_47[917]    = ( l_48 [472] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[918]    = ( l_48 [404] & !i[1699]) | ( l_48 [472] &  i[1699]);
assign l_47[919]    = ( l_48 [473] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[920]    = ( l_48 [404] & !i[1699]) | ( l_48 [473] &  i[1699]);
assign l_47[921]    = ( l_48 [474] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[922]    = ( l_48 [404] & !i[1699]) | ( l_48 [474] &  i[1699]);
assign l_47[923]    = ( l_48 [475] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[924]    = ( l_48 [404] & !i[1699]) | ( l_48 [475] &  i[1699]);
assign l_47[925]    = ( l_48 [476] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[926]    = ( l_48 [404] & !i[1699]) | ( l_48 [476] &  i[1699]);
assign l_47[927]    = ( l_48 [477] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[928]    = ( l_48 [404] & !i[1699]) | ( l_48 [477] &  i[1699]);
assign l_47[929]    = ( l_48 [478] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[930]    = ( l_48 [404] & !i[1699]) | ( l_48 [478] &  i[1699]);
assign l_47[931]    = ( l_48 [479] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[932]    = ( l_48 [404] & !i[1699]) | ( l_48 [479] &  i[1699]);
assign l_47[933]    = ( l_48 [480] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[934]    = ( l_48 [404] & !i[1699]) | ( l_48 [480] &  i[1699]);
assign l_47[935]    = ( l_48 [481] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[936]    = ( l_48 [404] & !i[1699]) | ( l_48 [481] &  i[1699]);
assign l_47[937]    = ( l_48 [482] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[938]    = ( l_48 [404] & !i[1699]) | ( l_48 [482] &  i[1699]);
assign l_47[939]    = ( l_48 [483] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[940]    = ( l_48 [404] & !i[1699]) | ( l_48 [483] &  i[1699]);
assign l_47[941]    = ( l_48 [484] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[942]    = ( l_48 [404] & !i[1699]) | ( l_48 [484] &  i[1699]);
assign l_47[943]    = ( l_48 [485] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[944]    = ( l_48 [404] & !i[1699]) | ( l_48 [485] &  i[1699]);
assign l_47[945]    = ( l_48 [486] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[946]    = ( l_48 [421] & !i[1699]) | ( l_48 [486] &  i[1699]);
assign l_47[947]    = ( l_48 [487] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[948]    = ( l_48 [421] & !i[1699]) | ( l_48 [487] &  i[1699]);
assign l_47[949]    = ( l_48 [488] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[950]    = ( l_48 [421] & !i[1699]) | ( l_48 [488] &  i[1699]);
assign l_47[951]    = ( l_48 [489] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[952]    = ( l_48 [421] & !i[1699]) | ( l_48 [489] &  i[1699]);
assign l_47[953]    = ( l_48 [490] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[954]    = ( l_48 [421] & !i[1699]) | ( l_48 [490] &  i[1699]);
assign l_47[955]    = ( l_48 [491] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[956]    = ( l_48 [421] & !i[1699]) | ( l_48 [491] &  i[1699]);
assign l_47[957]    = ( l_48 [492] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[958]    = ( l_48 [421] & !i[1699]) | ( l_48 [492] &  i[1699]);
assign l_47[959]    = ( l_48 [493] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[960]    = ( l_48 [421] & !i[1699]) | ( l_48 [493] &  i[1699]);
assign l_47[961]    = ( l_48 [494] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[962]    = ( l_48 [421] & !i[1699]) | ( l_48 [494] &  i[1699]);
assign l_47[963]    = ( l_48 [495] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[964]    = ( l_48 [421] & !i[1699]) | ( l_48 [495] &  i[1699]);
assign l_47[965]    = ( l_48 [496] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[966]    = ( l_48 [421] & !i[1699]) | ( l_48 [496] &  i[1699]);
assign l_47[967]    = ( l_48 [497] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[968]    = ( l_48 [421] & !i[1699]) | ( l_48 [497] &  i[1699]);
assign l_47[969]    = ( l_48 [498] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[970]    = ( l_48 [421] & !i[1699]) | ( l_48 [498] &  i[1699]);
assign l_47[971]    = ( l_48 [499] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[972]    = ( l_48 [421] & !i[1699]) | ( l_48 [499] &  i[1699]);
assign l_47[973]    = ( l_48 [500] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[974]    = ( l_48 [421] & !i[1699]) | ( l_48 [500] &  i[1699]);
assign l_47[975]    = ( l_48 [501] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[976]    = ( l_48 [421] & !i[1699]) | ( l_48 [501] &  i[1699]);
assign l_47[977]    = ( l_48 [502] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[978]    = ( l_48 [438] & !i[1699]) | ( l_48 [502] &  i[1699]);
assign l_47[979]    = ( l_48 [503] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[980]    = ( l_48 [438] & !i[1699]) | ( l_48 [503] &  i[1699]);
assign l_47[981]    = ( l_48 [504] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[982]    = ( l_48 [438] & !i[1699]) | ( l_48 [504] &  i[1699]);
assign l_47[983]    = ( l_48 [505] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[984]    = ( l_48 [438] & !i[1699]) | ( l_48 [505] &  i[1699]);
assign l_47[985]    = ( l_48 [506] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[986]    = ( l_48 [438] & !i[1699]) | ( l_48 [506] &  i[1699]);
assign l_47[987]    = ( l_48 [507] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[988]    = ( l_48 [438] & !i[1699]) | ( l_48 [507] &  i[1699]);
assign l_47[989]    = ( l_48 [508] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[990]    = ( l_48 [438] & !i[1699]) | ( l_48 [508] &  i[1699]);
assign l_47[991]    = ( l_48 [509] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[992]    = ( l_48 [438] & !i[1699]) | ( l_48 [509] &  i[1699]);
assign l_47[993]    = ( l_48 [510] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[994]    = ( l_48 [438] & !i[1699]) | ( l_48 [510] &  i[1699]);
assign l_47[995]    = ( l_48 [511] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[996]    = ( l_48 [438] & !i[1699]) | ( l_48 [511] &  i[1699]);
assign l_47[997]    = ( l_48 [512] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[998]    = ( l_48 [438] & !i[1699]) | ( l_48 [512] &  i[1699]);
assign l_47[999]    = ( l_48 [513] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[1000]    = ( l_48 [438] & !i[1699]) | ( l_48 [513] &  i[1699]);
assign l_47[1001]    = ( l_48 [514] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[1002]    = ( l_48 [438] & !i[1699]) | ( l_48 [514] &  i[1699]);
assign l_47[1003]    = ( l_48 [515] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[1004]    = ( l_48 [438] & !i[1699]) | ( l_48 [515] &  i[1699]);
assign l_47[1005]    = ( l_48 [516] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[1006]    = ( l_48 [438] & !i[1699]) | ( l_48 [516] &  i[1699]);
assign l_47[1007]    = ( l_48 [517] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[1008]    = ( l_48 [438] & !i[1699]) | ( l_48 [517] &  i[1699]);
assign l_47[1009]    = ( l_48 [518] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1010]    = ( l_48 [518] &  i[1699]);
assign l_47[1011]    = ( l_48 [519] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1012]    = ( l_48 [519] &  i[1699]);
assign l_47[1013]    = ( l_48 [520] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1014]    = ( l_48 [520] &  i[1699]);
assign l_47[1015]    = ( l_48 [521] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1016]    = ( l_48 [521] &  i[1699]);
assign l_47[1017]    = ( l_48 [522] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1018]    = ( l_48 [522] &  i[1699]);
assign l_47[1019]    = ( l_48 [523] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1020]    = ( l_48 [523] &  i[1699]);
assign l_47[1021]    = ( l_48 [524] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1022]    = ( l_48 [524] &  i[1699]);
assign l_47[1023]    = ( l_48 [525] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1024]    = ( l_48 [525] &  i[1699]);
assign l_47[1025]    = ( l_48 [526] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1026]    = ( l_48 [526] &  i[1699]);
assign l_47[1027]    = ( l_48 [527] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1028]    = ( l_48 [527] &  i[1699]);
assign l_47[1029]    = ( l_48 [528] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1030]    = ( l_48 [528] &  i[1699]);
assign l_47[1031]    = ( l_48 [529] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1032]    = ( l_48 [529] &  i[1699]);
assign l_47[1033]    = ( l_48 [530] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1034]    = ( l_48 [530] &  i[1699]);
assign l_47[1035]    = ( l_48 [531] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1036]    = ( l_48 [531] &  i[1699]);
assign l_47[1037]    = ( l_48 [532] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1038]    = ( l_48 [532] &  i[1699]);
assign l_47[1039]    = ( l_48 [533] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1040]    = ( l_48 [533] &  i[1699]);
assign l_47[1041]    = ( l_48 [534] & !i[1699]) | (      i[1699]);
assign l_47[1042]    = ( l_48 [272] & !i[1699]) | ( l_48 [534] &  i[1699]);
assign l_47[1043]    = ( l_48 [535] & !i[1699]) | ( l_48 [272] &  i[1699]);
assign l_47[1044]    = ( l_48 [289] & !i[1699]) | ( l_48 [535] &  i[1699]);
assign l_47[1045]    = ( l_48 [536] & !i[1699]) | ( l_48 [289] &  i[1699]);
assign l_47[1046]    = ( l_48 [306] & !i[1699]) | ( l_48 [536] &  i[1699]);
assign l_47[1047]    = ( l_48 [537] & !i[1699]) | ( l_48 [306] &  i[1699]);
assign l_47[1048]    = ( l_48 [338] & !i[1699]) | ( l_48 [537] &  i[1699]);
assign l_47[1049]    = ( l_48 [538] & !i[1699]) | ( l_48 [338] &  i[1699]);
assign l_47[1050]    = ( l_48 [404] & !i[1699]) | ( l_48 [538] &  i[1699]);
assign l_47[1051]    = ( l_48 [539] & !i[1699]) | ( l_48 [404] &  i[1699]);
assign l_47[1052]    = ( l_48 [421] & !i[1699]) | ( l_48 [539] &  i[1699]);
assign l_47[1053]    = ( l_48 [540] & !i[1699]) | ( l_48 [421] &  i[1699]);
assign l_47[1054]    = ( l_48 [438] & !i[1699]) | ( l_48 [540] &  i[1699]);
assign l_47[1055]    = ( l_48 [541] & !i[1699]) | ( l_48 [438] &  i[1699]);
assign l_47[1056]    = ( l_48 [541] &  i[1699]);
assign l_47[1057]    = ( l_48 [542]);
assign l_47[1058]    = ( l_48 [543]);
assign l_47[1059]    = ( l_48 [544]);
assign l_47[1060]    = ( l_48 [545]);
assign l_47[1061]    = ( l_48 [546]);
assign l_47[1062]    = ( l_48 [547]);
assign l_47[1063]    = ( l_48 [548]);
assign l_48[0]    = ( l_49 [0] & !i[1696]);
assign l_48[1]    = !i[1696];
assign l_48[2]    = ( l_49 [1] & !i[1696]);
assign l_48[3]    = ( l_49 [2] & !i[1696]);
assign l_48[4]    = ( l_49 [3] & !i[1696]);
assign l_48[5]    = ( l_49 [4] & !i[1696]);
assign l_48[6]    = ( l_49 [5] & !i[1696]);
assign l_48[7]    = ( l_49 [6] & !i[1696]);
assign l_48[8]    = ( l_49 [7] & !i[1696]);
assign l_48[9]    = ( l_49 [8] & !i[1696]);
assign l_48[10]    = ( l_49 [9] & !i[1696]);
assign l_48[11]    = ( l_49 [10] & !i[1696]);
assign l_48[12]    = ( l_49 [11] & !i[1696]);
assign l_48[13]    = ( l_49 [12] & !i[1696]);
assign l_48[14]    = ( l_49 [13] & !i[1696]);
assign l_48[15]    = ( l_49 [14] & !i[1696]);
assign l_48[16]    = ( l_49 [15] & !i[1696]);
assign l_48[17]    = ( l_49 [16] & !i[1696]);
assign l_48[18]    = ( l_49 [17] & !i[1696]);
assign l_48[19]    = ( l_49 [18] & !i[1696]);
assign l_48[20]    = ( l_49 [19] & !i[1696]);
assign l_48[21]    = ( l_49 [20] & !i[1696]);
assign l_48[22]    = ( l_49 [21] & !i[1696]);
assign l_48[23]    = ( l_49 [22] & !i[1696]);
assign l_48[24]    = ( l_49 [23] & !i[1696]);
assign l_48[25]    = ( l_49 [24] & !i[1696]);
assign l_48[26]    = ( l_49 [25] & !i[1696]);
assign l_48[27]    = ( l_49 [26] & !i[1696]);
assign l_48[28]    = ( l_49 [27] & !i[1696]);
assign l_48[29]    = ( l_49 [28] & !i[1696]);
assign l_48[30]    = ( l_49 [29] & !i[1696]);
assign l_48[31]    = ( l_49 [30] & !i[1696]);
assign l_48[32]    = ( l_49 [31] & !i[1696]);
assign l_48[33]    = ( l_49 [32] & !i[1696]);
assign l_48[34]    = ( l_49 [33] & !i[1696]);
assign l_48[35]    = ( l_49 [34] & !i[1696]);
assign l_48[36]    = ( l_49 [35] & !i[1696]);
assign l_48[37]    = ( l_49 [36] & !i[1696]);
assign l_48[38]    = ( l_49 [37] & !i[1696]);
assign l_48[39]    = ( l_49 [38] & !i[1696]);
assign l_48[40]    = ( l_49 [39] & !i[1696]);
assign l_48[41]    = ( l_49 [40] & !i[1696]);
assign l_48[42]    = ( l_49 [41] & !i[1696]);
assign l_48[43]    = ( l_49 [42] & !i[1696]);
assign l_48[44]    = ( l_49 [43] & !i[1696]);
assign l_48[45]    = ( l_49 [44] & !i[1696]);
assign l_48[46]    = ( l_49 [45] & !i[1696]);
assign l_48[47]    = ( l_49 [46] & !i[1696]);
assign l_48[48]    = ( l_49 [47] & !i[1696]);
assign l_48[49]    = ( l_49 [48] & !i[1696]);
assign l_48[50]    = ( l_49 [49] & !i[1696]);
assign l_48[51]    = ( l_49 [50] & !i[1696]);
assign l_48[52]    = ( l_49 [51] & !i[1696]);
assign l_48[53]    = ( l_49 [52] & !i[1696]);
assign l_48[54]    = ( l_49 [53] & !i[1696]);
assign l_48[55]    = ( l_49 [54] & !i[1696]);
assign l_48[56]    = ( l_49 [55] & !i[1696]);
assign l_48[57]    = ( l_49 [56] & !i[1696]);
assign l_48[58]    = ( l_49 [57] & !i[1696]);
assign l_48[59]    = ( l_49 [58] & !i[1696]);
assign l_48[60]    = ( l_49 [59] & !i[1696]);
assign l_48[61]    = ( l_49 [60] & !i[1696]);
assign l_48[62]    = ( l_49 [61] & !i[1696]);
assign l_48[63]    = ( l_49 [62] & !i[1696]);
assign l_48[64]    = ( l_49 [63] & !i[1696]);
assign l_48[65]    = ( l_49 [64] & !i[1696]);
assign l_48[66]    = ( l_49 [65] & !i[1696]);
assign l_48[67]    = ( l_49 [66] & !i[1696]);
assign l_48[68]    = ( l_49 [67] & !i[1696]);
assign l_48[69]    = ( l_49 [68] & !i[1696]);
assign l_48[70]    = ( l_49 [69] & !i[1696]);
assign l_48[71]    = ( l_49 [70] & !i[1696]);
assign l_48[72]    = ( l_49 [71] & !i[1696]);
assign l_48[73]    = ( l_49 [72] & !i[1696]);
assign l_48[74]    = ( l_49 [73] & !i[1696]);
assign l_48[75]    = ( l_49 [74] & !i[1696]);
assign l_48[76]    = ( l_49 [75] & !i[1696]);
assign l_48[77]    = ( l_49 [76] & !i[1696]);
assign l_48[78]    = ( l_49 [77] & !i[1696]);
assign l_48[79]    = ( l_49 [78] & !i[1696]);
assign l_48[80]    = ( l_49 [79] & !i[1696]);
assign l_48[81]    = ( l_49 [80] & !i[1696]);
assign l_48[82]    = ( l_49 [81] & !i[1696]);
assign l_48[83]    = ( l_49 [82] & !i[1696]);
assign l_48[84]    = ( l_49 [83] & !i[1696]);
assign l_48[85]    = ( l_49 [84] & !i[1696]);
assign l_48[86]    = ( l_49 [85] & !i[1696]);
assign l_48[87]    = ( l_49 [86] & !i[1696]);
assign l_48[88]    = ( l_49 [87] & !i[1696]);
assign l_48[89]    = ( l_49 [88] & !i[1696]);
assign l_48[90]    = ( l_49 [89] & !i[1696]);
assign l_48[91]    = ( l_49 [90] & !i[1696]);
assign l_48[92]    = ( l_49 [91] & !i[1696]);
assign l_48[93]    = ( l_49 [92] & !i[1696]);
assign l_48[94]    = ( l_49 [93] & !i[1696]);
assign l_48[95]    = ( l_49 [94] & !i[1696]);
assign l_48[96]    = ( l_49 [95] & !i[1696]);
assign l_48[97]    = ( l_49 [96] & !i[1696]);
assign l_48[98]    = ( l_49 [97] & !i[1696]);
assign l_48[99]    = ( l_49 [98] & !i[1696]);
assign l_48[100]    = ( l_49 [99] & !i[1696]);
assign l_48[101]    = ( l_49 [100] & !i[1696]);
assign l_48[102]    = ( l_49 [101] & !i[1696]);
assign l_48[103]    = ( l_49 [102] & !i[1696]);
assign l_48[104]    = ( l_49 [103] & !i[1696]);
assign l_48[105]    = ( l_49 [104] & !i[1696]);
assign l_48[106]    = ( l_49 [105] & !i[1696]);
assign l_48[107]    = ( l_49 [106] & !i[1696]);
assign l_48[108]    = ( l_49 [107] & !i[1696]);
assign l_48[109]    = ( l_49 [108] & !i[1696]);
assign l_48[110]    = ( l_49 [109] & !i[1696]);
assign l_48[111]    = ( l_49 [110] & !i[1696]);
assign l_48[112]    = ( l_49 [111] & !i[1696]);
assign l_48[113]    = ( l_49 [112] & !i[1696]);
assign l_48[114]    = ( l_49 [113] & !i[1696]);
assign l_48[115]    = ( l_49 [114] & !i[1696]);
assign l_48[116]    = ( l_49 [115] & !i[1696]);
assign l_48[117]    = ( l_49 [116] & !i[1696]);
assign l_48[118]    = ( l_49 [117] & !i[1696]);
assign l_48[119]    = ( l_49 [118] & !i[1696]);
assign l_48[120]    = ( l_49 [119] & !i[1696]);
assign l_48[121]    = ( l_49 [120] & !i[1696]);
assign l_48[122]    = ( l_49 [121] & !i[1696]);
assign l_48[123]    = ( l_49 [122] & !i[1696]);
assign l_48[124]    = ( l_49 [123] & !i[1696]);
assign l_48[125]    = ( l_49 [124] & !i[1696]);
assign l_48[126]    = ( l_49 [125] & !i[1696]);
assign l_48[127]    = ( l_49 [126] & !i[1696]);
assign l_48[128]    = ( l_49 [127] & !i[1696]);
assign l_48[129]    = ( l_49 [128] & !i[1696]);
assign l_48[130]    = ( l_49 [129] & !i[1696]);
assign l_48[131]    = ( l_49 [130] & !i[1696]);
assign l_48[132]    = (!i[1696]) | ( l_49 [0] &  i[1696]);
assign l_48[133]    = (!i[1696]) | ( l_49 [1] &  i[1696]);
assign l_48[134]    = (!i[1696]) | ( l_49 [2] &  i[1696]);
assign l_48[135]    = (!i[1696]) | ( l_49 [3] &  i[1696]);
assign l_48[136]    = (!i[1696]) | ( l_49 [4] &  i[1696]);
assign l_48[137]    = (!i[1696]) | ( l_49 [5] &  i[1696]);
assign l_48[138]    = (!i[1696]) | ( l_49 [6] &  i[1696]);
assign l_48[139]    = (!i[1696]) | ( l_49 [7] &  i[1696]);
assign l_48[140]    = (!i[1696]) | ( l_49 [8] &  i[1696]);
assign l_48[141]    = (!i[1696]) | ( l_49 [9] &  i[1696]);
assign l_48[142]    = (!i[1696]) | ( l_49 [10] &  i[1696]);
assign l_48[143]    = (!i[1696]) | ( l_49 [11] &  i[1696]);
assign l_48[144]    = (!i[1696]) | ( l_49 [12] &  i[1696]);
assign l_48[145]    = (!i[1696]) | ( l_49 [13] &  i[1696]);
assign l_48[146]    = (!i[1696]) | ( l_49 [14] &  i[1696]);
assign l_48[147]    = (!i[1696]) | ( l_49 [15] &  i[1696]);
assign l_48[148]    = (!i[1696]) | ( l_49 [16] &  i[1696]);
assign l_48[149]    = (!i[1696]) | ( l_49 [17] &  i[1696]);
assign l_48[150]    = (!i[1696]) | ( l_49 [18] &  i[1696]);
assign l_48[151]    = (!i[1696]) | ( l_49 [19] &  i[1696]);
assign l_48[152]    = (!i[1696]) | ( l_49 [20] &  i[1696]);
assign l_48[153]    = (!i[1696]) | ( l_49 [21] &  i[1696]);
assign l_48[154]    = (!i[1696]) | ( l_49 [22] &  i[1696]);
assign l_48[155]    = (!i[1696]) | ( l_49 [23] &  i[1696]);
assign l_48[156]    = (!i[1696]) | ( l_49 [24] &  i[1696]);
assign l_48[157]    = (!i[1696]) | ( l_49 [25] &  i[1696]);
assign l_48[158]    = (!i[1696]) | ( l_49 [26] &  i[1696]);
assign l_48[159]    = (!i[1696]) | ( l_49 [27] &  i[1696]);
assign l_48[160]    = (!i[1696]) | ( l_49 [28] &  i[1696]);
assign l_48[161]    = (!i[1696]) | ( l_49 [29] &  i[1696]);
assign l_48[162]    = (!i[1696]) | ( l_49 [30] &  i[1696]);
assign l_48[163]    = (!i[1696]) | ( l_49 [31] &  i[1696]);
assign l_48[164]    = (!i[1696]) | ( l_49 [32] &  i[1696]);
assign l_48[165]    = (!i[1696]) | ( l_49 [33] &  i[1696]);
assign l_48[166]    = (!i[1696]) | ( l_49 [34] &  i[1696]);
assign l_48[167]    = (!i[1696]) | ( l_49 [35] &  i[1696]);
assign l_48[168]    = (!i[1696]) | ( l_49 [36] &  i[1696]);
assign l_48[169]    = (!i[1696]) | ( l_49 [37] &  i[1696]);
assign l_48[170]    = (!i[1696]) | ( l_49 [38] &  i[1696]);
assign l_48[171]    = (!i[1696]) | ( l_49 [39] &  i[1696]);
assign l_48[172]    = (!i[1696]) | ( l_49 [40] &  i[1696]);
assign l_48[173]    = (!i[1696]) | ( l_49 [41] &  i[1696]);
assign l_48[174]    = (!i[1696]) | ( l_49 [42] &  i[1696]);
assign l_48[175]    = (!i[1696]) | ( l_49 [43] &  i[1696]);
assign l_48[176]    = (!i[1696]) | ( l_49 [44] &  i[1696]);
assign l_48[177]    = (!i[1696]) | ( l_49 [45] &  i[1696]);
assign l_48[178]    = (!i[1696]) | ( l_49 [46] &  i[1696]);
assign l_48[179]    = (!i[1696]) | ( l_49 [47] &  i[1696]);
assign l_48[180]    = (!i[1696]) | ( l_49 [48] &  i[1696]);
assign l_48[181]    = (!i[1696]) | ( l_49 [49] &  i[1696]);
assign l_48[182]    = (!i[1696]) | ( l_49 [50] &  i[1696]);
assign l_48[183]    = (!i[1696]) | ( l_49 [51] &  i[1696]);
assign l_48[184]    = (!i[1696]) | ( l_49 [52] &  i[1696]);
assign l_48[185]    = (!i[1696]) | ( l_49 [53] &  i[1696]);
assign l_48[186]    = (!i[1696]) | ( l_49 [54] &  i[1696]);
assign l_48[187]    = (!i[1696]) | ( l_49 [55] &  i[1696]);
assign l_48[188]    = (!i[1696]) | ( l_49 [56] &  i[1696]);
assign l_48[189]    = (!i[1696]) | ( l_49 [57] &  i[1696]);
assign l_48[190]    = (!i[1696]) | ( l_49 [58] &  i[1696]);
assign l_48[191]    = (!i[1696]) | ( l_49 [59] &  i[1696]);
assign l_48[192]    = (!i[1696]) | ( l_49 [60] &  i[1696]);
assign l_48[193]    = (!i[1696]) | ( l_49 [61] &  i[1696]);
assign l_48[194]    = (!i[1696]) | ( l_49 [62] &  i[1696]);
assign l_48[195]    = (!i[1696]) | ( l_49 [63] &  i[1696]);
assign l_48[196]    = (!i[1696]) | ( l_49 [64] &  i[1696]);
assign l_48[197]    = (!i[1696]) | ( l_49 [65] &  i[1696]);
assign l_48[198]    = (!i[1696]) | ( l_49 [66] &  i[1696]);
assign l_48[199]    = (!i[1696]) | ( l_49 [67] &  i[1696]);
assign l_48[200]    = (!i[1696]) | ( l_49 [68] &  i[1696]);
assign l_48[201]    = (!i[1696]) | ( l_49 [69] &  i[1696]);
assign l_48[202]    = (!i[1696]) | ( l_49 [70] &  i[1696]);
assign l_48[203]    = (!i[1696]) | ( l_49 [71] &  i[1696]);
assign l_48[204]    = (!i[1696]) | ( l_49 [72] &  i[1696]);
assign l_48[205]    = (!i[1696]) | ( l_49 [73] &  i[1696]);
assign l_48[206]    = (!i[1696]) | ( l_49 [74] &  i[1696]);
assign l_48[207]    = (!i[1696]) | ( l_49 [75] &  i[1696]);
assign l_48[208]    = (!i[1696]) | ( l_49 [76] &  i[1696]);
assign l_48[209]    = (!i[1696]) | ( l_49 [77] &  i[1696]);
assign l_48[210]    = (!i[1696]) | ( l_49 [78] &  i[1696]);
assign l_48[211]    = (!i[1696]) | ( l_49 [79] &  i[1696]);
assign l_48[212]    = (!i[1696]) | ( l_49 [80] &  i[1696]);
assign l_48[213]    = (!i[1696]) | ( l_49 [81] &  i[1696]);
assign l_48[214]    = (!i[1696]) | ( l_49 [82] &  i[1696]);
assign l_48[215]    = (!i[1696]) | ( l_49 [83] &  i[1696]);
assign l_48[216]    = (!i[1696]) | ( l_49 [84] &  i[1696]);
assign l_48[217]    = (!i[1696]) | ( l_49 [85] &  i[1696]);
assign l_48[218]    = (!i[1696]) | ( l_49 [86] &  i[1696]);
assign l_48[219]    = (!i[1696]) | ( l_49 [87] &  i[1696]);
assign l_48[220]    = (!i[1696]) | ( l_49 [88] &  i[1696]);
assign l_48[221]    = (!i[1696]) | ( l_49 [89] &  i[1696]);
assign l_48[222]    = (!i[1696]) | ( l_49 [90] &  i[1696]);
assign l_48[223]    = (!i[1696]) | ( l_49 [91] &  i[1696]);
assign l_48[224]    = (!i[1696]) | ( l_49 [92] &  i[1696]);
assign l_48[225]    = (!i[1696]) | ( l_49 [93] &  i[1696]);
assign l_48[226]    = (!i[1696]) | ( l_49 [94] &  i[1696]);
assign l_48[227]    = (!i[1696]) | ( l_49 [95] &  i[1696]);
assign l_48[228]    = (!i[1696]) | ( l_49 [96] &  i[1696]);
assign l_48[229]    = (!i[1696]) | ( l_49 [97] &  i[1696]);
assign l_48[230]    = (!i[1696]) | ( l_49 [98] &  i[1696]);
assign l_48[231]    = (!i[1696]) | ( l_49 [99] &  i[1696]);
assign l_48[232]    = (!i[1696]) | ( l_49 [100] &  i[1696]);
assign l_48[233]    = (!i[1696]) | ( l_49 [101] &  i[1696]);
assign l_48[234]    = (!i[1696]) | ( l_49 [102] &  i[1696]);
assign l_48[235]    = (!i[1696]) | ( l_49 [103] &  i[1696]);
assign l_48[236]    = (!i[1696]) | ( l_49 [104] &  i[1696]);
assign l_48[237]    = (!i[1696]) | ( l_49 [105] &  i[1696]);
assign l_48[238]    = (!i[1696]) | ( l_49 [106] &  i[1696]);
assign l_48[239]    = (!i[1696]) | ( l_49 [107] &  i[1696]);
assign l_48[240]    = (!i[1696]) | ( l_49 [108] &  i[1696]);
assign l_48[241]    = (!i[1696]) | ( l_49 [109] &  i[1696]);
assign l_48[242]    = (!i[1696]) | ( l_49 [110] &  i[1696]);
assign l_48[243]    = (!i[1696]) | ( l_49 [111] &  i[1696]);
assign l_48[244]    = (!i[1696]) | ( l_49 [112] &  i[1696]);
assign l_48[245]    = (!i[1696]) | ( l_49 [113] &  i[1696]);
assign l_48[246]    = (!i[1696]) | ( l_49 [114] &  i[1696]);
assign l_48[247]    = (!i[1696]) | ( l_49 [115] &  i[1696]);
assign l_48[248]    = (!i[1696]) | ( l_49 [116] &  i[1696]);
assign l_48[249]    = (!i[1696]) | ( l_49 [117] &  i[1696]);
assign l_48[250]    = (!i[1696]) | ( l_49 [118] &  i[1696]);
assign l_48[251]    = (!i[1696]) | ( l_49 [119] &  i[1696]);
assign l_48[252]    = (!i[1696]) | ( l_49 [120] &  i[1696]);
assign l_48[253]    = (!i[1696]) | ( l_49 [121] &  i[1696]);
assign l_48[254]    = (!i[1696]) | ( l_49 [122] &  i[1696]);
assign l_48[255]    = (!i[1696]) | ( l_49 [123] &  i[1696]);
assign l_48[256]    = (!i[1696]) | ( l_49 [124] &  i[1696]);
assign l_48[257]    = (!i[1696]) | ( l_49 [125] &  i[1696]);
assign l_48[258]    = (!i[1696]) | ( l_49 [126] &  i[1696]);
assign l_48[259]    = (!i[1696]) | ( l_49 [127] &  i[1696]);
assign l_48[260]    = (!i[1696]) | ( l_49 [128] &  i[1696]);
assign l_48[261]    = (!i[1696]) | ( l_49 [129] &  i[1696]);
assign l_48[262]    = (!i[1696]) | ( l_49 [130] &  i[1696]);
assign l_48[263]    = ( l_49 [131] & !i[1696]);
assign l_48[264]    = ( l_49 [132] & !i[1696]);
assign l_48[265]    = ( l_49 [133] & !i[1696]);
assign l_48[266]    = ( l_49 [134] & !i[1696]);
assign l_48[267]    = (!i[1696]) | ( l_49 [131] &  i[1696]);
assign l_48[268]    = (!i[1696]) | ( l_49 [132] &  i[1696]);
assign l_48[269]    = (!i[1696]) | ( l_49 [133] &  i[1696]);
assign l_48[270]    = (!i[1696]) | ( l_49 [134] &  i[1696]);
assign l_48[271]    = ( l_49 [0] & !i[1696]) | (      i[1696]);
assign l_48[272]    = ( l_49 [1] & !i[1696]) | (      i[1696]);
assign l_48[273]    = ( l_49 [2] & !i[1696]) | (      i[1696]);
assign l_48[274]    = ( l_49 [3] & !i[1696]) | (      i[1696]);
assign l_48[275]    = ( l_49 [4] & !i[1696]) | (      i[1696]);
assign l_48[276]    = ( l_49 [5] & !i[1696]) | (      i[1696]);
assign l_48[277]    = ( l_49 [6] & !i[1696]) | (      i[1696]);
assign l_48[278]    = ( l_49 [7] & !i[1696]) | (      i[1696]);
assign l_48[279]    = ( l_49 [8] & !i[1696]) | (      i[1696]);
assign l_48[280]    = ( l_49 [9] & !i[1696]) | (      i[1696]);
assign l_48[281]    = ( l_49 [10] & !i[1696]) | (      i[1696]);
assign l_48[282]    = ( l_49 [11] & !i[1696]) | (      i[1696]);
assign l_48[283]    = ( l_49 [12] & !i[1696]) | (      i[1696]);
assign l_48[284]    = ( l_49 [13] & !i[1696]) | (      i[1696]);
assign l_48[285]    = ( l_49 [14] & !i[1696]) | (      i[1696]);
assign l_48[286]    = ( l_49 [15] & !i[1696]) | (      i[1696]);
assign l_48[287]    = ( l_49 [16] & !i[1696]) | (      i[1696]);
assign l_48[288]    = ( l_49 [17] & !i[1696]) | (      i[1696]);
assign l_48[289]    = ( l_49 [18] & !i[1696]) | (      i[1696]);
assign l_48[290]    = ( l_49 [19] & !i[1696]) | (      i[1696]);
assign l_48[291]    = ( l_49 [20] & !i[1696]) | (      i[1696]);
assign l_48[292]    = ( l_49 [21] & !i[1696]) | (      i[1696]);
assign l_48[293]    = ( l_49 [22] & !i[1696]) | (      i[1696]);
assign l_48[294]    = ( l_49 [23] & !i[1696]) | (      i[1696]);
assign l_48[295]    = ( l_49 [24] & !i[1696]) | (      i[1696]);
assign l_48[296]    = ( l_49 [25] & !i[1696]) | (      i[1696]);
assign l_48[297]    = ( l_49 [26] & !i[1696]) | (      i[1696]);
assign l_48[298]    = ( l_49 [27] & !i[1696]) | (      i[1696]);
assign l_48[299]    = ( l_49 [28] & !i[1696]) | (      i[1696]);
assign l_48[300]    = ( l_49 [29] & !i[1696]) | (      i[1696]);
assign l_48[301]    = ( l_49 [30] & !i[1696]) | (      i[1696]);
assign l_48[302]    = ( l_49 [31] & !i[1696]) | (      i[1696]);
assign l_48[303]    = ( l_49 [32] & !i[1696]) | (      i[1696]);
assign l_48[304]    = ( l_49 [33] & !i[1696]) | (      i[1696]);
assign l_48[305]    = ( l_49 [34] & !i[1696]) | (      i[1696]);
assign l_48[306]    = ( l_49 [35] & !i[1696]) | (      i[1696]);
assign l_48[307]    = ( l_49 [36] & !i[1696]) | (      i[1696]);
assign l_48[308]    = ( l_49 [37] & !i[1696]) | (      i[1696]);
assign l_48[309]    = ( l_49 [38] & !i[1696]) | (      i[1696]);
assign l_48[310]    = ( l_49 [39] & !i[1696]) | (      i[1696]);
assign l_48[311]    = ( l_49 [40] & !i[1696]) | (      i[1696]);
assign l_48[312]    = ( l_49 [41] & !i[1696]) | (      i[1696]);
assign l_48[313]    = ( l_49 [42] & !i[1696]) | (      i[1696]);
assign l_48[314]    = ( l_49 [43] & !i[1696]) | (      i[1696]);
assign l_48[315]    = ( l_49 [44] & !i[1696]) | (      i[1696]);
assign l_48[316]    = ( l_49 [45] & !i[1696]) | (      i[1696]);
assign l_48[317]    = ( l_49 [46] & !i[1696]) | (      i[1696]);
assign l_48[318]    = ( l_49 [47] & !i[1696]) | (      i[1696]);
assign l_48[319]    = ( l_49 [48] & !i[1696]) | (      i[1696]);
assign l_48[320]    = ( l_49 [49] & !i[1696]) | (      i[1696]);
assign l_48[321]    = ( l_49 [50] & !i[1696]) | (      i[1696]);
assign l_48[322]    = ( l_49 [51] & !i[1696]) | (      i[1696]);
assign l_48[323]    = ( l_49 [52] & !i[1696]) | (      i[1696]);
assign l_48[324]    = ( l_49 [53] & !i[1696]) | (      i[1696]);
assign l_48[325]    = ( l_49 [54] & !i[1696]) | (      i[1696]);
assign l_48[326]    = ( l_49 [55] & !i[1696]) | (      i[1696]);
assign l_48[327]    = ( l_49 [56] & !i[1696]) | (      i[1696]);
assign l_48[328]    = ( l_49 [57] & !i[1696]) | (      i[1696]);
assign l_48[329]    = ( l_49 [58] & !i[1696]) | (      i[1696]);
assign l_48[330]    = ( l_49 [59] & !i[1696]) | (      i[1696]);
assign l_48[331]    = ( l_49 [60] & !i[1696]) | (      i[1696]);
assign l_48[332]    = ( l_49 [61] & !i[1696]) | (      i[1696]);
assign l_48[333]    = ( l_49 [62] & !i[1696]) | (      i[1696]);
assign l_48[334]    = ( l_49 [63] & !i[1696]) | (      i[1696]);
assign l_48[335]    = ( l_49 [64] & !i[1696]) | (      i[1696]);
assign l_48[336]    = ( l_49 [65] & !i[1696]) | (      i[1696]);
assign l_48[337]    = ( l_49 [66] & !i[1696]) | (      i[1696]);
assign l_48[338]    =  i[1696];
assign l_48[339]    = ( l_49 [67] & !i[1696]) | (      i[1696]);
assign l_48[340]    = ( l_49 [68] & !i[1696]) | (      i[1696]);
assign l_48[341]    = ( l_49 [69] & !i[1696]) | (      i[1696]);
assign l_48[342]    = ( l_49 [70] & !i[1696]) | (      i[1696]);
assign l_48[343]    = ( l_49 [71] & !i[1696]) | (      i[1696]);
assign l_48[344]    = ( l_49 [72] & !i[1696]) | (      i[1696]);
assign l_48[345]    = ( l_49 [73] & !i[1696]) | (      i[1696]);
assign l_48[346]    = ( l_49 [74] & !i[1696]) | (      i[1696]);
assign l_48[347]    = ( l_49 [75] & !i[1696]) | (      i[1696]);
assign l_48[348]    = ( l_49 [76] & !i[1696]) | (      i[1696]);
assign l_48[349]    = ( l_49 [77] & !i[1696]) | (      i[1696]);
assign l_48[350]    = ( l_49 [78] & !i[1696]) | (      i[1696]);
assign l_48[351]    = ( l_49 [79] & !i[1696]) | (      i[1696]);
assign l_48[352]    = ( l_49 [80] & !i[1696]) | (      i[1696]);
assign l_48[353]    = ( l_49 [81] & !i[1696]) | (      i[1696]);
assign l_48[354]    = ( l_49 [82] & !i[1696]) | (      i[1696]);
assign l_48[355]    = ( l_49 [83] & !i[1696]) | (      i[1696]);
assign l_48[356]    = ( l_49 [84] & !i[1696]) | (      i[1696]);
assign l_48[357]    = ( l_49 [85] & !i[1696]) | (      i[1696]);
assign l_48[358]    = ( l_49 [86] & !i[1696]) | (      i[1696]);
assign l_48[359]    = ( l_49 [87] & !i[1696]) | (      i[1696]);
assign l_48[360]    = ( l_49 [88] & !i[1696]) | (      i[1696]);
assign l_48[361]    = ( l_49 [89] & !i[1696]) | (      i[1696]);
assign l_48[362]    = ( l_49 [90] & !i[1696]) | (      i[1696]);
assign l_48[363]    = ( l_49 [91] & !i[1696]) | (      i[1696]);
assign l_48[364]    = ( l_49 [92] & !i[1696]) | (      i[1696]);
assign l_48[365]    = ( l_49 [93] & !i[1696]) | (      i[1696]);
assign l_48[366]    = ( l_49 [94] & !i[1696]) | (      i[1696]);
assign l_48[367]    = ( l_49 [95] & !i[1696]) | (      i[1696]);
assign l_48[368]    = ( l_49 [96] & !i[1696]) | (      i[1696]);
assign l_48[369]    = ( l_49 [97] & !i[1696]) | (      i[1696]);
assign l_48[370]    = ( l_49 [98] & !i[1696]) | (      i[1696]);
assign l_48[371]    = ( l_49 [99] & !i[1696]) | (      i[1696]);
assign l_48[372]    = ( l_49 [100] & !i[1696]) | (      i[1696]);
assign l_48[373]    = ( l_49 [101] & !i[1696]) | (      i[1696]);
assign l_48[374]    = ( l_49 [102] & !i[1696]) | (      i[1696]);
assign l_48[375]    = ( l_49 [103] & !i[1696]) | (      i[1696]);
assign l_48[376]    = ( l_49 [104] & !i[1696]) | (      i[1696]);
assign l_48[377]    = ( l_49 [105] & !i[1696]) | (      i[1696]);
assign l_48[378]    = ( l_49 [106] & !i[1696]) | (      i[1696]);
assign l_48[379]    = ( l_49 [107] & !i[1696]) | (      i[1696]);
assign l_48[380]    = ( l_49 [108] & !i[1696]) | (      i[1696]);
assign l_48[381]    = ( l_49 [109] & !i[1696]) | (      i[1696]);
assign l_48[382]    = ( l_49 [110] & !i[1696]) | (      i[1696]);
assign l_48[383]    = ( l_49 [111] & !i[1696]) | (      i[1696]);
assign l_48[384]    = ( l_49 [112] & !i[1696]) | (      i[1696]);
assign l_48[385]    = ( l_49 [113] & !i[1696]) | (      i[1696]);
assign l_48[386]    = ( l_49 [114] & !i[1696]) | (      i[1696]);
assign l_48[387]    = ( l_49 [115] & !i[1696]) | (      i[1696]);
assign l_48[388]    = ( l_49 [116] & !i[1696]) | (      i[1696]);
assign l_48[389]    = ( l_49 [117] & !i[1696]) | (      i[1696]);
assign l_48[390]    = ( l_49 [118] & !i[1696]) | (      i[1696]);
assign l_48[391]    = ( l_49 [119] & !i[1696]) | (      i[1696]);
assign l_48[392]    = ( l_49 [120] & !i[1696]) | (      i[1696]);
assign l_48[393]    = ( l_49 [121] & !i[1696]) | (      i[1696]);
assign l_48[394]    = ( l_49 [122] & !i[1696]) | (      i[1696]);
assign l_48[395]    = ( l_49 [123] & !i[1696]) | (      i[1696]);
assign l_48[396]    = ( l_49 [124] & !i[1696]) | (      i[1696]);
assign l_48[397]    = ( l_49 [125] & !i[1696]) | (      i[1696]);
assign l_48[398]    = ( l_49 [126] & !i[1696]) | (      i[1696]);
assign l_48[399]    = ( l_49 [127] & !i[1696]) | (      i[1696]);
assign l_48[400]    = ( l_49 [128] & !i[1696]) | (      i[1696]);
assign l_48[401]    = ( l_49 [129] & !i[1696]) | (      i[1696]);
assign l_48[402]    = ( l_49 [130] & !i[1696]) | (      i[1696]);
assign l_48[403]    = ( l_49 [0] &  i[1696]);
assign l_48[404]    = ( l_49 [1] &  i[1696]);
assign l_48[405]    = ( l_49 [2] &  i[1696]);
assign l_48[406]    = ( l_49 [3] &  i[1696]);
assign l_48[407]    = ( l_49 [4] &  i[1696]);
assign l_48[408]    = ( l_49 [5] &  i[1696]);
assign l_48[409]    = ( l_49 [6] &  i[1696]);
assign l_48[410]    = ( l_49 [7] &  i[1696]);
assign l_48[411]    = ( l_49 [8] &  i[1696]);
assign l_48[412]    = ( l_49 [9] &  i[1696]);
assign l_48[413]    = ( l_49 [10] &  i[1696]);
assign l_48[414]    = ( l_49 [11] &  i[1696]);
assign l_48[415]    = ( l_49 [12] &  i[1696]);
assign l_48[416]    = ( l_49 [13] &  i[1696]);
assign l_48[417]    = ( l_49 [14] &  i[1696]);
assign l_48[418]    = ( l_49 [15] &  i[1696]);
assign l_48[419]    = ( l_49 [16] &  i[1696]);
assign l_48[420]    = ( l_49 [17] &  i[1696]);
assign l_48[421]    = ( l_49 [18] &  i[1696]);
assign l_48[422]    = ( l_49 [19] &  i[1696]);
assign l_48[423]    = ( l_49 [20] &  i[1696]);
assign l_48[424]    = ( l_49 [21] &  i[1696]);
assign l_48[425]    = ( l_49 [22] &  i[1696]);
assign l_48[426]    = ( l_49 [23] &  i[1696]);
assign l_48[427]    = ( l_49 [24] &  i[1696]);
assign l_48[428]    = ( l_49 [25] &  i[1696]);
assign l_48[429]    = ( l_49 [26] &  i[1696]);
assign l_48[430]    = ( l_49 [27] &  i[1696]);
assign l_48[431]    = ( l_49 [28] &  i[1696]);
assign l_48[432]    = ( l_49 [29] &  i[1696]);
assign l_48[433]    = ( l_49 [30] &  i[1696]);
assign l_48[434]    = ( l_49 [31] &  i[1696]);
assign l_48[435]    = ( l_49 [32] &  i[1696]);
assign l_48[436]    = ( l_49 [33] &  i[1696]);
assign l_48[437]    = ( l_49 [34] &  i[1696]);
assign l_48[438]    = ( l_49 [35] &  i[1696]);
assign l_48[439]    = ( l_49 [36] &  i[1696]);
assign l_48[440]    = ( l_49 [37] &  i[1696]);
assign l_48[441]    = ( l_49 [38] &  i[1696]);
assign l_48[442]    = ( l_49 [39] &  i[1696]);
assign l_48[443]    = ( l_49 [40] &  i[1696]);
assign l_48[444]    = ( l_49 [41] &  i[1696]);
assign l_48[445]    = ( l_49 [42] &  i[1696]);
assign l_48[446]    = ( l_49 [43] &  i[1696]);
assign l_48[447]    = ( l_49 [44] &  i[1696]);
assign l_48[448]    = ( l_49 [45] &  i[1696]);
assign l_48[449]    = ( l_49 [46] &  i[1696]);
assign l_48[450]    = ( l_49 [47] &  i[1696]);
assign l_48[451]    = ( l_49 [48] &  i[1696]);
assign l_48[452]    = ( l_49 [49] &  i[1696]);
assign l_48[453]    = ( l_49 [50] &  i[1696]);
assign l_48[454]    = ( l_49 [51] &  i[1696]);
assign l_48[455]    = ( l_49 [52] &  i[1696]);
assign l_48[456]    = ( l_49 [53] &  i[1696]);
assign l_48[457]    = ( l_49 [54] &  i[1696]);
assign l_48[458]    = ( l_49 [55] &  i[1696]);
assign l_48[459]    = ( l_49 [56] &  i[1696]);
assign l_48[460]    = ( l_49 [57] &  i[1696]);
assign l_48[461]    = ( l_49 [58] &  i[1696]);
assign l_48[462]    = ( l_49 [59] &  i[1696]);
assign l_48[463]    = ( l_49 [60] &  i[1696]);
assign l_48[464]    = ( l_49 [61] &  i[1696]);
assign l_48[465]    = ( l_49 [62] &  i[1696]);
assign l_48[466]    = ( l_49 [63] &  i[1696]);
assign l_48[467]    = ( l_49 [64] &  i[1696]);
assign l_48[468]    = ( l_49 [65] &  i[1696]);
assign l_48[469]    = ( l_49 [66] &  i[1696]);
assign l_48[470]    = ( l_49 [67] &  i[1696]);
assign l_48[471]    = ( l_49 [68] &  i[1696]);
assign l_48[472]    = ( l_49 [69] &  i[1696]);
assign l_48[473]    = ( l_49 [70] &  i[1696]);
assign l_48[474]    = ( l_49 [71] &  i[1696]);
assign l_48[475]    = ( l_49 [72] &  i[1696]);
assign l_48[476]    = ( l_49 [73] &  i[1696]);
assign l_48[477]    = ( l_49 [74] &  i[1696]);
assign l_48[478]    = ( l_49 [75] &  i[1696]);
assign l_48[479]    = ( l_49 [76] &  i[1696]);
assign l_48[480]    = ( l_49 [77] &  i[1696]);
assign l_48[481]    = ( l_49 [78] &  i[1696]);
assign l_48[482]    = ( l_49 [79] &  i[1696]);
assign l_48[483]    = ( l_49 [80] &  i[1696]);
assign l_48[484]    = ( l_49 [81] &  i[1696]);
assign l_48[485]    = ( l_49 [82] &  i[1696]);
assign l_48[486]    = ( l_49 [83] &  i[1696]);
assign l_48[487]    = ( l_49 [84] &  i[1696]);
assign l_48[488]    = ( l_49 [85] &  i[1696]);
assign l_48[489]    = ( l_49 [86] &  i[1696]);
assign l_48[490]    = ( l_49 [87] &  i[1696]);
assign l_48[491]    = ( l_49 [88] &  i[1696]);
assign l_48[492]    = ( l_49 [89] &  i[1696]);
assign l_48[493]    = ( l_49 [90] &  i[1696]);
assign l_48[494]    = ( l_49 [91] &  i[1696]);
assign l_48[495]    = ( l_49 [92] &  i[1696]);
assign l_48[496]    = ( l_49 [93] &  i[1696]);
assign l_48[497]    = ( l_49 [94] &  i[1696]);
assign l_48[498]    = ( l_49 [95] &  i[1696]);
assign l_48[499]    = ( l_49 [96] &  i[1696]);
assign l_48[500]    = ( l_49 [97] &  i[1696]);
assign l_48[501]    = ( l_49 [98] &  i[1696]);
assign l_48[502]    = ( l_49 [99] &  i[1696]);
assign l_48[503]    = ( l_49 [100] &  i[1696]);
assign l_48[504]    = ( l_49 [101] &  i[1696]);
assign l_48[505]    = ( l_49 [102] &  i[1696]);
assign l_48[506]    = ( l_49 [103] &  i[1696]);
assign l_48[507]    = ( l_49 [104] &  i[1696]);
assign l_48[508]    = ( l_49 [105] &  i[1696]);
assign l_48[509]    = ( l_49 [106] &  i[1696]);
assign l_48[510]    = ( l_49 [107] &  i[1696]);
assign l_48[511]    = ( l_49 [108] &  i[1696]);
assign l_48[512]    = ( l_49 [109] &  i[1696]);
assign l_48[513]    = ( l_49 [110] &  i[1696]);
assign l_48[514]    = ( l_49 [111] &  i[1696]);
assign l_48[515]    = ( l_49 [112] &  i[1696]);
assign l_48[516]    = ( l_49 [113] &  i[1696]);
assign l_48[517]    = ( l_49 [114] &  i[1696]);
assign l_48[518]    = ( l_49 [115] &  i[1696]);
assign l_48[519]    = ( l_49 [116] &  i[1696]);
assign l_48[520]    = ( l_49 [117] &  i[1696]);
assign l_48[521]    = ( l_49 [118] &  i[1696]);
assign l_48[522]    = ( l_49 [119] &  i[1696]);
assign l_48[523]    = ( l_49 [120] &  i[1696]);
assign l_48[524]    = ( l_49 [121] &  i[1696]);
assign l_48[525]    = ( l_49 [122] &  i[1696]);
assign l_48[526]    = ( l_49 [123] &  i[1696]);
assign l_48[527]    = ( l_49 [124] &  i[1696]);
assign l_48[528]    = ( l_49 [125] &  i[1696]);
assign l_48[529]    = ( l_49 [126] &  i[1696]);
assign l_48[530]    = ( l_49 [127] &  i[1696]);
assign l_48[531]    = ( l_49 [128] &  i[1696]);
assign l_48[532]    = ( l_49 [129] &  i[1696]);
assign l_48[533]    = ( l_49 [130] &  i[1696]);
assign l_48[534]    = ( l_49 [131] & !i[1696]) | (      i[1696]);
assign l_48[535]    = ( l_49 [132] & !i[1696]) | (      i[1696]);
assign l_48[536]    = ( l_49 [133] & !i[1696]) | (      i[1696]);
assign l_48[537]    = ( l_49 [134] & !i[1696]) | (      i[1696]);
assign l_48[538]    = ( l_49 [131] &  i[1696]);
assign l_48[539]    = ( l_49 [132] &  i[1696]);
assign l_48[540]    = ( l_49 [133] &  i[1696]);
assign l_48[541]    = ( l_49 [134] &  i[1696]);
assign l_48[542]    = ( l_49 [135]);
assign l_48[543]    = ( l_49 [136]);
assign l_48[544]    = ( l_49 [137]);
assign l_48[545]    = ( l_49 [138]);
assign l_48[546]    = ( l_49 [139]);
assign l_48[547]    = ( l_49 [140]);
assign l_48[548]    = ( l_49 [141]);
assign l_49[0]    = ( l_50 [0]);
assign l_49[1]    = ( l_50 [1]);
assign l_49[2]    = ( l_50 [2] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[3]    = ( l_50 [3] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[4]    = ( l_50 [4] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[5]    = ( l_50 [5] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[6]    = ( l_50 [6] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[7]    = ( l_50 [7] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[8]    = ( l_50 [8] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[9]    = ( l_50 [9] & !i[1825]) | ( l_50 [0] &  i[1825]);
assign l_49[10]    = ( l_50 [9] & !i[1825]) | ( l_50 [2] &  i[1825]);
assign l_49[11]    = ( l_50 [9] & !i[1825]) | ( l_50 [3] &  i[1825]);
assign l_49[12]    = ( l_50 [9] & !i[1825]) | ( l_50 [4] &  i[1825]);
assign l_49[13]    = ( l_50 [9] & !i[1825]) | ( l_50 [5] &  i[1825]);
assign l_49[14]    = ( l_50 [9] & !i[1825]) | ( l_50 [6] &  i[1825]);
assign l_49[15]    = ( l_50 [9] & !i[1825]) | ( l_50 [7] &  i[1825]);
assign l_49[16]    = ( l_50 [9] & !i[1825]) | ( l_50 [8] &  i[1825]);
assign l_49[17]    = ( l_50 [10]);
assign l_49[18]    = ( l_50 [11]);
assign l_49[19]    = ( l_50 [12] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[20]    = ( l_50 [13] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[21]    = ( l_50 [14] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[22]    = ( l_50 [15] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[23]    = ( l_50 [16] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[24]    = ( l_50 [17] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[25]    = ( l_50 [18] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[26]    = ( l_50 [19] & !i[1825]) | ( l_50 [10] &  i[1825]);
assign l_49[27]    = ( l_50 [19] & !i[1825]) | ( l_50 [12] &  i[1825]);
assign l_49[28]    = ( l_50 [19] & !i[1825]) | ( l_50 [13] &  i[1825]);
assign l_49[29]    = ( l_50 [19] & !i[1825]) | ( l_50 [14] &  i[1825]);
assign l_49[30]    = ( l_50 [19] & !i[1825]) | ( l_50 [15] &  i[1825]);
assign l_49[31]    = ( l_50 [19] & !i[1825]) | ( l_50 [16] &  i[1825]);
assign l_49[32]    = ( l_50 [19] & !i[1825]) | ( l_50 [17] &  i[1825]);
assign l_49[33]    = ( l_50 [19] & !i[1825]) | ( l_50 [18] &  i[1825]);
assign l_49[34]    = ( l_50 [20]);
assign l_49[35]    = ( l_50 [21]);
assign l_49[36]    = ( l_50 [22] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[37]    = ( l_50 [23] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[38]    = ( l_50 [24] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[39]    = ( l_50 [25] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[40]    = ( l_50 [26] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[41]    = ( l_50 [27] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[42]    = ( l_50 [28] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[43]    = ( l_50 [29] & !i[1825]) | ( l_50 [20] &  i[1825]);
assign l_49[44]    = ( l_50 [29] & !i[1825]) | ( l_50 [22] &  i[1825]);
assign l_49[45]    = ( l_50 [29] & !i[1825]) | ( l_50 [23] &  i[1825]);
assign l_49[46]    = ( l_50 [29] & !i[1825]) | ( l_50 [24] &  i[1825]);
assign l_49[47]    = ( l_50 [29] & !i[1825]) | ( l_50 [25] &  i[1825]);
assign l_49[48]    = ( l_50 [29] & !i[1825]) | ( l_50 [26] &  i[1825]);
assign l_49[49]    = ( l_50 [29] & !i[1825]) | ( l_50 [27] &  i[1825]);
assign l_49[50]    = ( l_50 [29] & !i[1825]) | ( l_50 [28] &  i[1825]);
assign l_49[51]    = ( l_50 [30]);
assign l_49[52]    = ( l_50 [31] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[53]    = ( l_50 [32] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[54]    = ( l_50 [33] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[55]    = ( l_50 [34] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[56]    = ( l_50 [35] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[57]    = ( l_50 [36] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[58]    = ( l_50 [37] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[59]    = ( l_50 [38] & !i[1825]) | ( l_50 [30] &  i[1825]);
assign l_49[60]    = ( l_50 [38] & !i[1825]) | ( l_50 [31] &  i[1825]);
assign l_49[61]    = ( l_50 [38] & !i[1825]) | ( l_50 [32] &  i[1825]);
assign l_49[62]    = ( l_50 [38] & !i[1825]) | ( l_50 [33] &  i[1825]);
assign l_49[63]    = ( l_50 [38] & !i[1825]) | ( l_50 [34] &  i[1825]);
assign l_49[64]    = ( l_50 [38] & !i[1825]) | ( l_50 [35] &  i[1825]);
assign l_49[65]    = ( l_50 [38] & !i[1825]) | ( l_50 [36] &  i[1825]);
assign l_49[66]    = ( l_50 [38] & !i[1825]) | ( l_50 [37] &  i[1825]);
assign l_49[67]    = ( l_50 [9]);
assign l_49[68]    = ( l_50 [39] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[69]    = ( l_50 [40] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[70]    = ( l_50 [41] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[71]    = ( l_50 [42] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[72]    = ( l_50 [43] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[73]    = ( l_50 [44] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[74]    = ( l_50 [45] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[75]    = ( l_50 [46] & !i[1825]) | ( l_50 [9] &  i[1825]);
assign l_49[76]    = ( l_50 [46] & !i[1825]) | ( l_50 [39] &  i[1825]);
assign l_49[77]    = ( l_50 [46] & !i[1825]) | ( l_50 [40] &  i[1825]);
assign l_49[78]    = ( l_50 [46] & !i[1825]) | ( l_50 [41] &  i[1825]);
assign l_49[79]    = ( l_50 [46] & !i[1825]) | ( l_50 [42] &  i[1825]);
assign l_49[80]    = ( l_50 [46] & !i[1825]) | ( l_50 [43] &  i[1825]);
assign l_49[81]    = ( l_50 [46] & !i[1825]) | ( l_50 [44] &  i[1825]);
assign l_49[82]    = ( l_50 [46] & !i[1825]) | ( l_50 [45] &  i[1825]);
assign l_49[83]    = ( l_50 [19]);
assign l_49[84]    = ( l_50 [47] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[85]    = ( l_50 [48] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[86]    = ( l_50 [49] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[87]    = ( l_50 [50] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[88]    = ( l_50 [51] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[89]    = ( l_50 [52] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[90]    = ( l_50 [53] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[91]    = ( l_50 [54] & !i[1825]) | ( l_50 [19] &  i[1825]);
assign l_49[92]    = ( l_50 [54] & !i[1825]) | ( l_50 [47] &  i[1825]);
assign l_49[93]    = ( l_50 [54] & !i[1825]) | ( l_50 [48] &  i[1825]);
assign l_49[94]    = ( l_50 [54] & !i[1825]) | ( l_50 [49] &  i[1825]);
assign l_49[95]    = ( l_50 [54] & !i[1825]) | ( l_50 [50] &  i[1825]);
assign l_49[96]    = ( l_50 [54] & !i[1825]) | ( l_50 [51] &  i[1825]);
assign l_49[97]    = ( l_50 [54] & !i[1825]) | ( l_50 [52] &  i[1825]);
assign l_49[98]    = ( l_50 [54] & !i[1825]) | ( l_50 [53] &  i[1825]);
assign l_49[99]    = ( l_50 [29]);
assign l_49[100]    = ( l_50 [55] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[101]    = ( l_50 [56] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[102]    = ( l_50 [57] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[103]    = ( l_50 [58] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[104]    = ( l_50 [59] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[105]    = ( l_50 [60] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[106]    = ( l_50 [61] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[107]    = ( l_50 [62] & !i[1825]) | ( l_50 [29] &  i[1825]);
assign l_49[108]    = ( l_50 [62] & !i[1825]) | ( l_50 [55] &  i[1825]);
assign l_49[109]    = ( l_50 [62] & !i[1825]) | ( l_50 [56] &  i[1825]);
assign l_49[110]    = ( l_50 [62] & !i[1825]) | ( l_50 [57] &  i[1825]);
assign l_49[111]    = ( l_50 [62] & !i[1825]) | ( l_50 [58] &  i[1825]);
assign l_49[112]    = ( l_50 [62] & !i[1825]) | ( l_50 [59] &  i[1825]);
assign l_49[113]    = ( l_50 [62] & !i[1825]) | ( l_50 [60] &  i[1825]);
assign l_49[114]    = ( l_50 [62] & !i[1825]) | ( l_50 [61] &  i[1825]);
assign l_49[115]    = ( l_50 [38]);
assign l_49[116]    = ( l_50 [63] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[117]    = ( l_50 [64] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[118]    = ( l_50 [65] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[119]    = ( l_50 [66] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[120]    = ( l_50 [67] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[121]    = ( l_50 [68] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[122]    = ( l_50 [69] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[123]    = ( l_50 [70] & !i[1825]) | ( l_50 [38] &  i[1825]);
assign l_49[124]    = ( l_50 [70] & !i[1825]) | ( l_50 [63] &  i[1825]);
assign l_49[125]    = ( l_50 [70] & !i[1825]) | ( l_50 [64] &  i[1825]);
assign l_49[126]    = ( l_50 [70] & !i[1825]) | ( l_50 [65] &  i[1825]);
assign l_49[127]    = ( l_50 [70] & !i[1825]) | ( l_50 [66] &  i[1825]);
assign l_49[128]    = ( l_50 [70] & !i[1825]) | ( l_50 [67] &  i[1825]);
assign l_49[129]    = ( l_50 [70] & !i[1825]) | ( l_50 [68] &  i[1825]);
assign l_49[130]    = ( l_50 [70] & !i[1825]) | ( l_50 [69] &  i[1825]);
assign l_49[131]    = ( l_50 [46]);
assign l_49[132]    = ( l_50 [54]);
assign l_49[133]    = ( l_50 [62]);
assign l_49[134]    = ( l_50 [70]);
assign l_49[135]    =  i[1825];
assign l_49[136]    = ( l_50 [71]);
assign l_49[137]    = ( l_50 [72]);
assign l_49[138]    = ( l_50 [73]);
assign l_49[139]    = ( l_50 [74]);
assign l_49[140]    = ( l_50 [75]);
assign l_49[141]    = ( l_50 [76]);
assign l_50[0]    = ( l_51 [0]);
assign l_50[1]    = ( l_51 [1]);
assign l_50[2]    = ( l_51 [2] & !i[1827]) | ( l_51 [0] &  i[1827]);
assign l_50[3]    = ( l_51 [3] & !i[1827]) | ( l_51 [0] &  i[1827]);
assign l_50[4]    = ( l_51 [2] & !i[1827]) | ( l_51 [3] &  i[1827]);
assign l_50[5]    = ( l_51 [2]);
assign l_50[6]    = ( l_51 [4] & !i[1827]) | ( l_51 [2] &  i[1827]);
assign l_50[7]    = ( l_51 [5] & !i[1827]) | ( l_51 [2] &  i[1827]);
assign l_50[8]    = ( l_51 [4] & !i[1827]) | ( l_51 [5] &  i[1827]);
assign l_50[9]    = ( l_51 [4]);
assign l_50[10]    = ( l_51 [6]);
assign l_50[11]    = ( l_51 [7]);
assign l_50[12]    = ( l_51 [8] & !i[1827]) | ( l_51 [6] &  i[1827]);
assign l_50[13]    = ( l_51 [9] & !i[1827]) | ( l_51 [6] &  i[1827]);
assign l_50[14]    = ( l_51 [8] & !i[1827]) | ( l_51 [9] &  i[1827]);
assign l_50[15]    = ( l_51 [8]);
assign l_50[16]    = ( l_51 [10] & !i[1827]) | ( l_51 [8] &  i[1827]);
assign l_50[17]    = ( l_51 [11] & !i[1827]) | ( l_51 [8] &  i[1827]);
assign l_50[18]    = ( l_51 [10] & !i[1827]) | ( l_51 [11] &  i[1827]);
assign l_50[19]    = ( l_51 [10]);
assign l_50[20]    = ( l_51 [12]);
assign l_50[21]    = ( l_51 [13]);
assign l_50[22]    = ( l_51 [14] & !i[1827]) | ( l_51 [12] &  i[1827]);
assign l_50[23]    = ( l_51 [15] & !i[1827]) | ( l_51 [12] &  i[1827]);
assign l_50[24]    = ( l_51 [14] & !i[1827]) | ( l_51 [15] &  i[1827]);
assign l_50[25]    = ( l_51 [14]);
assign l_50[26]    = ( l_51 [16] & !i[1827]) | ( l_51 [14] &  i[1827]);
assign l_50[27]    = ( l_51 [17] & !i[1827]) | ( l_51 [14] &  i[1827]);
assign l_50[28]    = ( l_51 [16] & !i[1827]) | ( l_51 [17] &  i[1827]);
assign l_50[29]    = ( l_51 [16]);
assign l_50[30]    = ( l_51 [18]);
assign l_50[31]    = ( l_51 [19] & !i[1827]) | ( l_51 [18] &  i[1827]);
assign l_50[32]    = ( l_51 [20] & !i[1827]) | ( l_51 [18] &  i[1827]);
assign l_50[33]    = ( l_51 [19] & !i[1827]) | ( l_51 [20] &  i[1827]);
assign l_50[34]    = ( l_51 [19]);
assign l_50[35]    = ( l_51 [21] & !i[1827]) | ( l_51 [19] &  i[1827]);
assign l_50[36]    = ( l_51 [22] & !i[1827]) | ( l_51 [19] &  i[1827]);
assign l_50[37]    = ( l_51 [21] & !i[1827]) | ( l_51 [22] &  i[1827]);
assign l_50[38]    = ( l_51 [21]);
assign l_50[39]    = ( l_51 [23] & !i[1827]) | ( l_51 [4] &  i[1827]);
assign l_50[40]    = ( l_51 [24] & !i[1827]) | ( l_51 [4] &  i[1827]);
assign l_50[41]    = ( l_51 [23] & !i[1827]) | ( l_51 [24] &  i[1827]);
assign l_50[42]    = ( l_51 [23]);
assign l_50[43]    = ( l_51 [25] & !i[1827]) | ( l_51 [23] &  i[1827]);
assign l_50[44]    = ( l_51 [26] & !i[1827]) | ( l_51 [23] &  i[1827]);
assign l_50[45]    = ( l_51 [25] & !i[1827]) | ( l_51 [26] &  i[1827]);
assign l_50[46]    = ( l_51 [25]);
assign l_50[47]    = ( l_51 [27] & !i[1827]) | ( l_51 [10] &  i[1827]);
assign l_50[48]    = ( l_51 [28] & !i[1827]) | ( l_51 [10] &  i[1827]);
assign l_50[49]    = ( l_51 [27] & !i[1827]) | ( l_51 [28] &  i[1827]);
assign l_50[50]    = ( l_51 [27]);
assign l_50[51]    = ( l_51 [29] & !i[1827]) | ( l_51 [27] &  i[1827]);
assign l_50[52]    = ( l_51 [30] & !i[1827]) | ( l_51 [27] &  i[1827]);
assign l_50[53]    = ( l_51 [29] & !i[1827]) | ( l_51 [30] &  i[1827]);
assign l_50[54]    = ( l_51 [29]);
assign l_50[55]    = ( l_51 [31] & !i[1827]) | ( l_51 [16] &  i[1827]);
assign l_50[56]    = ( l_51 [32] & !i[1827]) | ( l_51 [16] &  i[1827]);
assign l_50[57]    = ( l_51 [31] & !i[1827]) | ( l_51 [32] &  i[1827]);
assign l_50[58]    = ( l_51 [31]);
assign l_50[59]    = ( l_51 [33] & !i[1827]) | ( l_51 [31] &  i[1827]);
assign l_50[60]    = ( l_51 [34] & !i[1827]) | ( l_51 [31] &  i[1827]);
assign l_50[61]    = ( l_51 [33] & !i[1827]) | ( l_51 [34] &  i[1827]);
assign l_50[62]    = ( l_51 [33]);
assign l_50[63]    = ( l_51 [35] & !i[1827]) | ( l_51 [21] &  i[1827]);
assign l_50[64]    = ( l_51 [36] & !i[1827]) | ( l_51 [21] &  i[1827]);
assign l_50[65]    = ( l_51 [35] & !i[1827]) | ( l_51 [36] &  i[1827]);
assign l_50[66]    = ( l_51 [35]);
assign l_50[67]    = ( l_51 [37] & !i[1827]) | ( l_51 [35] &  i[1827]);
assign l_50[68]    = ( l_51 [38] & !i[1827]) | ( l_51 [35] &  i[1827]);
assign l_50[69]    = ( l_51 [37] & !i[1827]) | ( l_51 [38] &  i[1827]);
assign l_50[70]    = ( l_51 [37]);
assign l_50[71]    =  i[1827];
assign l_50[72]    = ( l_51 [39]);
assign l_50[73]    = ( l_51 [40]);
assign l_50[74]    = ( l_51 [41]);
assign l_50[75]    = ( l_51 [42]);
assign l_50[76]    = ( l_51 [43]);
assign l_51[0]    = ( l_52 [0] & !i[1823]) | ( l_52 [1] &  i[1823]);
assign l_51[1]    = ( l_52 [2]);
assign l_51[2]    = ( l_52 [3] & !i[1823]) | ( l_52 [4] &  i[1823]);
assign l_51[3]    = ( l_52 [5] & !i[1823]) | ( l_52 [6] &  i[1823]);
assign l_51[4]    = ( l_52 [7] & !i[1823]) | ( l_52 [8] &  i[1823]);
assign l_51[5]    = ( l_52 [9] & !i[1823]) | ( l_52 [10] &  i[1823]);
assign l_51[6]    = ( l_52 [11] & !i[1823]) | ( l_52 [12] &  i[1823]);
assign l_51[7]    = ( l_52 [13]);
assign l_51[8]    = ( l_52 [14] & !i[1823]) | ( l_52 [15] &  i[1823]);
assign l_51[9]    = ( l_52 [16] & !i[1823]) | ( l_52 [17] &  i[1823]);
assign l_51[10]    = ( l_52 [18] & !i[1823]) | ( l_52 [19] &  i[1823]);
assign l_51[11]    = ( l_52 [20] & !i[1823]) | ( l_52 [21] &  i[1823]);
assign l_51[12]    = ( l_52 [22] & !i[1823]) | ( l_52 [23] &  i[1823]);
assign l_51[13]    = ( l_52 [24]);
assign l_51[14]    = ( l_52 [25] & !i[1823]) | ( l_52 [26] &  i[1823]);
assign l_51[15]    = ( l_52 [27] & !i[1823]) | ( l_52 [28] &  i[1823]);
assign l_51[16]    = ( l_52 [29] & !i[1823]) | ( l_52 [30] &  i[1823]);
assign l_51[17]    = ( l_52 [31] & !i[1823]) | ( l_52 [32] &  i[1823]);
assign l_51[18]    = ( l_52 [33] & !i[1823]) | ( l_52 [34] &  i[1823]);
assign l_51[19]    = ( l_52 [35] & !i[1823]) | ( l_52 [36] &  i[1823]);
assign l_51[20]    = ( l_52 [37] & !i[1823]) | ( l_52 [38] &  i[1823]);
assign l_51[21]    = ( l_52 [39] & !i[1823]) | ( l_52 [40] &  i[1823]);
assign l_51[22]    = ( l_52 [41] & !i[1823]) | ( l_52 [42] &  i[1823]);
assign l_51[23]    = ( l_52 [43] & !i[1823]) | ( l_52 [44] &  i[1823]);
assign l_51[24]    = ( l_52 [45] & !i[1823]) | ( l_52 [46] &  i[1823]);
assign l_51[25]    = ( l_52 [47] & !i[1823]) | ( l_52 [0] &  i[1823]);
assign l_51[26]    = ( l_52 [48] & !i[1823]) | ( l_52 [49] &  i[1823]);
assign l_51[27]    = ( l_52 [50] & !i[1823]) | ( l_52 [51] &  i[1823]);
assign l_51[28]    = ( l_52 [52] & !i[1823]) | ( l_52 [53] &  i[1823]);
assign l_51[29]    = ( l_52 [54] & !i[1823]) | ( l_52 [11] &  i[1823]);
assign l_51[30]    = ( l_52 [55] & !i[1823]) | ( l_52 [56] &  i[1823]);
assign l_51[31]    = ( l_52 [57] & !i[1823]) | ( l_52 [58] &  i[1823]);
assign l_51[32]    = ( l_52 [59] & !i[1823]) | ( l_52 [60] &  i[1823]);
assign l_51[33]    = ( l_52 [61] & !i[1823]) | ( l_52 [22] &  i[1823]);
assign l_51[34]    = ( l_52 [62] & !i[1823]) | ( l_52 [63] &  i[1823]);
assign l_51[35]    = ( l_52 [64] & !i[1823]) | ( l_52 [65] &  i[1823]);
assign l_51[36]    = ( l_52 [66] & !i[1823]) | ( l_52 [67] &  i[1823]);
assign l_51[37]    = ( l_52 [68] & !i[1823]) | ( l_52 [33] &  i[1823]);
assign l_51[38]    = ( l_52 [69] & !i[1823]) | ( l_52 [70] &  i[1823]);
assign l_51[39]    =  i[1823];
assign l_51[40]    = ( l_52 [71]);
assign l_51[41]    = ( l_52 [72]);
assign l_51[42]    = ( l_52 [73]);
assign l_51[43]    = ( l_52 [74]);
assign l_52[0]    = ( l_53 [0]);
assign l_52[1]    = ( l_53 [1]);
assign l_52[2]    = ( l_53 [2]);
assign l_52[3]    = ( l_53 [3]);
assign l_52[4]    = ( l_53 [4]);
assign l_52[5]    = ( l_53 [3] & !i[1828]) | ( l_53 [0] &  i[1828]);
assign l_52[6]    = ( l_53 [4] & !i[1828]) | ( l_53 [1] &  i[1828]);
assign l_52[7]    = ( l_53 [5]);
assign l_52[8]    = ( l_53 [6]);
assign l_52[9]    = ( l_53 [5] & !i[1828]) | ( l_53 [3] &  i[1828]);
assign l_52[10]    = ( l_53 [6] & !i[1828]) | ( l_53 [4] &  i[1828]);
assign l_52[11]    = ( l_53 [7]);
assign l_52[12]    = ( l_53 [8]);
assign l_52[13]    = ( l_53 [9]);
assign l_52[14]    = ( l_53 [10]);
assign l_52[15]    = ( l_53 [11]);
assign l_52[16]    = ( l_53 [10] & !i[1828]) | ( l_53 [7] &  i[1828]);
assign l_52[17]    = ( l_53 [11] & !i[1828]) | ( l_53 [8] &  i[1828]);
assign l_52[18]    = ( l_53 [12]);
assign l_52[19]    = ( l_53 [13]);
assign l_52[20]    = ( l_53 [12] & !i[1828]) | ( l_53 [10] &  i[1828]);
assign l_52[21]    = ( l_53 [13] & !i[1828]) | ( l_53 [11] &  i[1828]);
assign l_52[22]    = ( l_53 [14]);
assign l_52[23]    = ( l_53 [15]);
assign l_52[24]    = ( l_53 [16]);
assign l_52[25]    = ( l_53 [17]);
assign l_52[26]    = ( l_53 [18]);
assign l_52[27]    = ( l_53 [17] & !i[1828]) | ( l_53 [14] &  i[1828]);
assign l_52[28]    = ( l_53 [18] & !i[1828]) | ( l_53 [15] &  i[1828]);
assign l_52[29]    = ( l_53 [19]);
assign l_52[30]    = ( l_53 [20]);
assign l_52[31]    = ( l_53 [19] & !i[1828]) | ( l_53 [17] &  i[1828]);
assign l_52[32]    = ( l_53 [20] & !i[1828]) | ( l_53 [18] &  i[1828]);
assign l_52[33]    = ( l_53 [21]);
assign l_52[34]    = ( l_53 [22]);
assign l_52[35]    = ( l_53 [23]);
assign l_52[36]    = ( l_53 [24]);
assign l_52[37]    = ( l_53 [23] & !i[1828]) | ( l_53 [21] &  i[1828]);
assign l_52[38]    = ( l_53 [24] & !i[1828]) | ( l_53 [22] &  i[1828]);
assign l_52[39]    = ( l_53 [25]);
assign l_52[40]    = ( l_53 [26]);
assign l_52[41]    = ( l_53 [25] & !i[1828]) | ( l_53 [23] &  i[1828]);
assign l_52[42]    = ( l_53 [26] & !i[1828]) | ( l_53 [24] &  i[1828]);
assign l_52[43]    = ( l_53 [27]);
assign l_52[44]    = ( l_53 [28]);
assign l_52[45]    = ( l_53 [27] & !i[1828]) | ( l_53 [5] &  i[1828]);
assign l_52[46]    = ( l_53 [28] & !i[1828]) | ( l_53 [6] &  i[1828]);
assign l_52[47]    = ( l_53 [29]);
assign l_52[48]    = ( l_53 [29] & !i[1828]) | ( l_53 [27] &  i[1828]);
assign l_52[49]    = ( l_53 [0] & !i[1828]) | ( l_53 [28] &  i[1828]);
assign l_52[50]    = ( l_53 [30]);
assign l_52[51]    = ( l_53 [31]);
assign l_52[52]    = ( l_53 [30] & !i[1828]) | ( l_53 [12] &  i[1828]);
assign l_52[53]    = ( l_53 [31] & !i[1828]) | ( l_53 [13] &  i[1828]);
assign l_52[54]    = ( l_53 [32]);
assign l_52[55]    = ( l_53 [32] & !i[1828]) | ( l_53 [30] &  i[1828]);
assign l_52[56]    = ( l_53 [7] & !i[1828]) | ( l_53 [31] &  i[1828]);
assign l_52[57]    = ( l_53 [33]);
assign l_52[58]    = ( l_53 [34]);
assign l_52[59]    = ( l_53 [33] & !i[1828]) | ( l_53 [19] &  i[1828]);
assign l_52[60]    = ( l_53 [34] & !i[1828]) | ( l_53 [20] &  i[1828]);
assign l_52[61]    = ( l_53 [35]);
assign l_52[62]    = ( l_53 [35] & !i[1828]) | ( l_53 [33] &  i[1828]);
assign l_52[63]    = ( l_53 [14] & !i[1828]) | ( l_53 [34] &  i[1828]);
assign l_52[64]    = ( l_53 [36]);
assign l_52[65]    = ( l_53 [37]);
assign l_52[66]    = ( l_53 [36] & !i[1828]) | ( l_53 [25] &  i[1828]);
assign l_52[67]    = ( l_53 [37] & !i[1828]) | ( l_53 [26] &  i[1828]);
assign l_52[68]    = ( l_53 [38]);
assign l_52[69]    = ( l_53 [38] & !i[1828]) | ( l_53 [36] &  i[1828]);
assign l_52[70]    = ( l_53 [21] & !i[1828]) | ( l_53 [37] &  i[1828]);
assign l_52[71]    =  i[1828];
assign l_52[72]    = ( l_53 [39]);
assign l_52[73]    = ( l_53 [40]);
assign l_52[74]    = ( l_53 [41]);
assign l_53[0]    = ( l_54 [0]);
assign l_53[1]    = ( l_54 [1]);
assign l_53[2]    = ( l_54 [2]);
assign l_53[3]    = ( l_54 [3] & !i[1824]) | ( l_54 [0] &  i[1824]);
assign l_53[4]    = ( l_54 [4] & !i[1824]) | ( l_54 [1] &  i[1824]);
assign l_53[5]    = ( l_54 [5] & !i[1824]) | ( l_54 [0] &  i[1824]);
assign l_53[6]    = ( l_54 [0] & !i[1824]) | ( l_54 [1] &  i[1824]);
assign l_53[7]    = ( l_54 [6]);
assign l_53[8]    = ( l_54 [7]);
assign l_53[9]    = ( l_54 [8]);
assign l_53[10]    = ( l_54 [9] & !i[1824]) | ( l_54 [6] &  i[1824]);
assign l_53[11]    = ( l_54 [10] & !i[1824]) | ( l_54 [7] &  i[1824]);
assign l_53[12]    = ( l_54 [11] & !i[1824]) | ( l_54 [6] &  i[1824]);
assign l_53[13]    = ( l_54 [6] & !i[1824]) | ( l_54 [7] &  i[1824]);
assign l_53[14]    = ( l_54 [12]);
assign l_53[15]    = ( l_54 [13]);
assign l_53[16]    = ( l_54 [14]);
assign l_53[17]    = ( l_54 [15] & !i[1824]) | ( l_54 [12] &  i[1824]);
assign l_53[18]    = ( l_54 [16] & !i[1824]) | ( l_54 [13] &  i[1824]);
assign l_53[19]    = ( l_54 [17] & !i[1824]) | ( l_54 [12] &  i[1824]);
assign l_53[20]    = ( l_54 [12] & !i[1824]) | ( l_54 [13] &  i[1824]);
assign l_53[21]    = ( l_54 [18]);
assign l_53[22]    = ( l_54 [19]);
assign l_53[23]    = ( l_54 [20] & !i[1824]) | ( l_54 [18] &  i[1824]);
assign l_53[24]    = ( l_54 [21] & !i[1824]) | ( l_54 [19] &  i[1824]);
assign l_53[25]    = ( l_54 [22] & !i[1824]) | ( l_54 [18] &  i[1824]);
assign l_53[26]    = ( l_54 [18] & !i[1824]) | ( l_54 [19] &  i[1824]);
assign l_53[27]    = ( l_54 [5] & !i[1824]) | ( l_54 [3] &  i[1824]);
assign l_53[28]    = ( l_54 [0] & !i[1824]) | ( l_54 [4] &  i[1824]);
assign l_53[29]    = ( l_54 [5]);
assign l_53[30]    = ( l_54 [11] & !i[1824]) | ( l_54 [9] &  i[1824]);
assign l_53[31]    = ( l_54 [6] & !i[1824]) | ( l_54 [10] &  i[1824]);
assign l_53[32]    = ( l_54 [11]);
assign l_53[33]    = ( l_54 [17] & !i[1824]) | ( l_54 [15] &  i[1824]);
assign l_53[34]    = ( l_54 [12] & !i[1824]) | ( l_54 [16] &  i[1824]);
assign l_53[35]    = ( l_54 [17]);
assign l_53[36]    = ( l_54 [22] & !i[1824]) | ( l_54 [20] &  i[1824]);
assign l_53[37]    = ( l_54 [18] & !i[1824]) | ( l_54 [21] &  i[1824]);
assign l_53[38]    = ( l_54 [22]);
assign l_53[39]    =  i[1824];
assign l_53[40]    = ( l_54 [23]);
assign l_53[41]    = ( l_54 [24]);
assign l_54[0]    = ( l_55 [0]);
assign l_54[1]    = ( l_55 [1]);
assign l_54[2]    = ( l_55 [2]);
assign l_54[3]    = ( l_55 [3] & !i[1826]) | ( l_55 [0] &  i[1826]);
assign l_54[4]    = ( l_55 [0] & !i[1826]) | ( l_55 [1] &  i[1826]);
assign l_54[5]    = ( l_55 [3]);
assign l_54[6]    = ( l_55 [4]);
assign l_54[7]    = ( l_55 [5]);
assign l_54[8]    = ( l_55 [6]);
assign l_54[9]    = ( l_55 [7] & !i[1826]) | ( l_55 [4] &  i[1826]);
assign l_54[10]    = ( l_55 [4] & !i[1826]) | ( l_55 [5] &  i[1826]);
assign l_54[11]    = ( l_55 [7]);
assign l_54[12]    = ( l_55 [8]);
assign l_54[13]    = ( l_55 [9]);
assign l_54[14]    = ( l_55 [10]);
assign l_54[15]    = ( l_55 [11] & !i[1826]) | ( l_55 [8] &  i[1826]);
assign l_54[16]    = ( l_55 [8] & !i[1826]) | ( l_55 [9] &  i[1826]);
assign l_54[17]    = ( l_55 [11]);
assign l_54[18]    = ( l_55 [12]);
assign l_54[19]    = ( l_55 [13]);
assign l_54[20]    = ( l_55 [14] & !i[1826]) | ( l_55 [12] &  i[1826]);
assign l_54[21]    = ( l_55 [12] & !i[1826]) | ( l_55 [13] &  i[1826]);
assign l_54[22]    = ( l_55 [14]);
assign l_54[23]    =  i[1826];
assign l_54[24]    = ( l_55 [15]);
assign l_55[0]    = ( l_56 [0] & !i[1822]) | ( l_56 [1] &  i[1822]);
assign l_55[1]    = ( l_56 [2] & !i[1822]) | ( l_56 [3] &  i[1822]);
assign l_55[2]    = ( l_56 [3]);
assign l_55[3]    = (!i[1822]) | ( l_56 [2] &  i[1822]);
assign l_55[4]    = ( l_56 [4] & !i[1822]) | ( l_56 [5] &  i[1822]);
assign l_55[5]    = ( l_56 [6] & !i[1822]) | ( l_56 [7] &  i[1822]);
assign l_55[6]    = ( l_56 [7]);
assign l_55[7]    = ( l_56 [3] & !i[1822]) | ( l_56 [6] &  i[1822]);
assign l_55[8]    = ( l_56 [8] & !i[1822]) | ( l_56 [9] &  i[1822]);
assign l_55[9]    = ( l_56 [10] & !i[1822]) | ( l_56 [11] &  i[1822]);
assign l_55[10]    = ( l_56 [11]);
assign l_55[11]    = ( l_56 [7] & !i[1822]) | ( l_56 [10] &  i[1822]);
assign l_55[12]    = ( l_56 [12] & !i[1822]) | ( l_56 [13] &  i[1822]);
assign l_55[13]    = ( l_56 [14] & !i[1822]);
assign l_55[14]    = ( l_56 [11] & !i[1822]) | ( l_56 [14] &  i[1822]);
assign l_55[15]    =  i[1822];
assign l_56[0]    = ( l_57 [0] & !i[1698]) | (      i[1698]);
assign l_56[1]    = ( l_57 [1] & !i[1698]) | (      i[1698]);
assign l_56[2]    = ( l_57 [2] & !i[1698]) | (      i[1698]);
assign l_56[3]    = ( l_57 [3] & !i[1698]) | (      i[1698]);
assign l_56[4]    = ( l_57 [3] & !i[1698]) | ( l_57 [0] &  i[1698]);
assign l_56[5]    = ( l_57 [3] & !i[1698]) | ( l_57 [1] &  i[1698]);
assign l_56[6]    = ( l_57 [3] & !i[1698]) | ( l_57 [2] &  i[1698]);
assign l_56[7]    = ( l_57 [3]);
assign l_56[8]    = ( l_57 [4] & !i[1698]) | ( l_57 [3] &  i[1698]);
assign l_56[9]    = ( l_57 [5] & !i[1698]) | ( l_57 [3] &  i[1698]);
assign l_56[10]    = ( l_57 [6] & !i[1698]) | ( l_57 [3] &  i[1698]);
assign l_56[11]    = ( l_57 [3] &  i[1698]);
assign l_56[12]    = ( l_57 [4] &  i[1698]);
assign l_56[13]    = ( l_57 [5] &  i[1698]);
assign l_56[14]    = ( l_57 [6] &  i[1698]);
assign l_57[0]    = ( l_58 [0] & !i[1701]) | (      i[1701]);
assign l_57[1]    = ( l_58 [1] & !i[1701]) | ( l_58 [0] &  i[1701]);
assign l_57[2]    = ( l_58 [0]);
assign l_57[3]    = ( l_58 [1]);
assign l_57[4]    = ( l_58 [2] & !i[1701]) | ( l_58 [1] &  i[1701]);
assign l_57[5]    = ( l_58 [2] &  i[1701]);
assign l_57[6]    = ( l_58 [2]);
assign l_58[0]    = ( l_59 [0] & !i[1700]) | (      i[1700]);
assign l_58[1]    = ( l_59 [0]);
assign l_58[2]    = ( l_59 [0] &  i[1700]);
assign l_59[0]    =  i[1697];

endmodule
