module module_output_bit_63(i,o);

input [1893:0] i;
output  o;

wire [0:0] l_0;
wire [1:0] l_1;
wire [3:0] l_2;
wire [7:0] l_3;
wire [13:0] l_4;
wire [13:0] l_5;
wire [13:0] l_6;
wire [13:0] l_7;
wire [19:0] l_8;
wire [17:0] l_9;
wire [17:0] l_10;
wire [17:0] l_11;
wire [17:0] l_12;
wire [17:0] l_13;
wire [17:0] l_14;
wire [17:0] l_15;
wire [17:0] l_16;
wire [12:0] l_17;
wire [12:0] l_18;
wire [18:0] l_19;
wire [23:0] l_20;

assign	l_20[23:0]	= 24'b0;

assign o = l_0[0];

assign l_0[0]    = ( l_1 [0] & !i[63]) | ( l_1 [1] &  i[63]);
assign l_1[0]    = ( l_2 [0] & !i[1713]) | ( l_2 [1] &  i[1713]);
assign l_1[1]    = ( l_2 [2] & !i[1713]) | ( l_2 [3] &  i[1713]);
assign l_2[0]    = ( l_3 [0] & !i[1714]) | ( l_3 [1] &  i[1714]);
assign l_2[1]    = ( l_3 [2] & !i[1714]) | ( l_3 [3] &  i[1714]);
assign l_2[2]    = ( l_3 [4] & !i[1714]) | ( l_3 [5] &  i[1714]);
assign l_2[3]    = ( l_3 [6] & !i[1714]) | ( l_3 [7] &  i[1714]);
assign l_3[0]    = ( l_4 [0] &  i[1715]);
assign l_3[1]    = ( l_4 [1] & !i[1715]) | ( l_4 [2] &  i[1715]);
assign l_3[2]    = ( l_4 [3] & !i[1715]) | ( l_4 [4] &  i[1715]);
assign l_3[3]    = ( l_4 [5] & !i[1715]) | ( l_4 [6] &  i[1715]);
assign l_3[4]    = (!i[1715]) | ( l_4 [7] &  i[1715]);
assign l_3[5]    = ( l_4 [8] & !i[1715]) | ( l_4 [9] &  i[1715]);
assign l_3[6]    = ( l_4 [10] & !i[1715]) | ( l_4 [11] &  i[1715]);
assign l_3[7]    = ( l_4 [12] & !i[1715]) | ( l_4 [13] &  i[1715]);
assign l_4[0]    = ( l_5 [0] & !i[1716]);
assign l_4[1]    = ( l_5 [1] & !i[1716]);
assign l_4[2]    = ( l_5 [2] & !i[1716]);
assign l_4[3]    = ( l_5 [3] & !i[1716]);
assign l_4[4]    = ( l_5 [4] & !i[1716]);
assign l_4[5]    = ( l_5 [5] & !i[1716]);
assign l_4[6]    = ( l_5 [6] & !i[1716]);
assign l_4[7]    = ( l_5 [7] & !i[1716]) | (      i[1716]);
assign l_4[8]    = ( l_5 [8] & !i[1716]) | (      i[1716]);
assign l_4[9]    = ( l_5 [9] & !i[1716]) | (      i[1716]);
assign l_4[10]    = ( l_5 [10] & !i[1716]) | (      i[1716]);
assign l_4[11]    = ( l_5 [11] & !i[1716]) | (      i[1716]);
assign l_4[12]    = ( l_5 [12] & !i[1716]) | (      i[1716]);
assign l_4[13]    = ( l_5 [13] & !i[1716]) | (      i[1716]);
assign l_5[0]    = ( l_6 [0] & !i[1717]);
assign l_5[1]    = ( l_6 [1] & !i[1717]);
assign l_5[2]    = ( l_6 [2] & !i[1717]);
assign l_5[3]    = ( l_6 [3] & !i[1717]);
assign l_5[4]    = ( l_6 [4] & !i[1717]);
assign l_5[5]    = ( l_6 [5] & !i[1717]);
assign l_5[6]    = ( l_6 [6] & !i[1717]);
assign l_5[7]    = ( l_6 [7] & !i[1717]) | (      i[1717]);
assign l_5[8]    = ( l_6 [8] & !i[1717]) | (      i[1717]);
assign l_5[9]    = ( l_6 [9] & !i[1717]) | (      i[1717]);
assign l_5[10]    = ( l_6 [10] & !i[1717]) | (      i[1717]);
assign l_5[11]    = ( l_6 [11] & !i[1717]) | (      i[1717]);
assign l_5[12]    = ( l_6 [12] & !i[1717]) | (      i[1717]);
assign l_5[13]    = ( l_6 [13] & !i[1717]) | (      i[1717]);
assign l_6[0]    = ( l_7 [0] &  i[1723]);
assign l_6[1]    = ( l_7 [1] &  i[1723]);
assign l_6[2]    = ( l_7 [2] &  i[1723]);
assign l_6[3]    = ( l_7 [3] &  i[1723]);
assign l_6[4]    = ( l_7 [4] &  i[1723]);
assign l_6[5]    = ( l_7 [5] &  i[1723]);
assign l_6[6]    = ( l_7 [6] &  i[1723]);
assign l_6[7]    = (!i[1723]) | ( l_7 [7] &  i[1723]);
assign l_6[8]    = (!i[1723]) | ( l_7 [8] &  i[1723]);
assign l_6[9]    = (!i[1723]) | ( l_7 [9] &  i[1723]);
assign l_6[10]    = (!i[1723]) | ( l_7 [10] &  i[1723]);
assign l_6[11]    = (!i[1723]) | ( l_7 [11] &  i[1723]);
assign l_6[12]    = (!i[1723]) | ( l_7 [12] &  i[1723]);
assign l_6[13]    = (!i[1723]) | ( l_7 [13] &  i[1723]);
assign l_7[0]    = ( l_8 [0] & !i[1707]);
assign l_7[1]    = ( l_8 [1] & !i[1707]) | ( l_8 [2] &  i[1707]);
assign l_7[2]    = ( l_8 [3] & !i[1707]) | ( l_8 [4] &  i[1707]);
assign l_7[3]    = ( l_8 [5] & !i[1707]) | ( l_8 [6] &  i[1707]);
assign l_7[4]    = ( l_8 [7] & !i[1707]) | ( l_8 [8] &  i[1707]);
assign l_7[5]    = ( l_8 [5] & !i[1707]) | ( l_8 [9] &  i[1707]);
assign l_7[6]    = ( l_8 [5] &  i[1707]);
assign l_7[7]    = ( l_8 [10] & !i[1707]) | ( l_8 [11] &  i[1707]);
assign l_7[8]    = ( l_8 [12] & !i[1707]) | ( l_8 [13] &  i[1707]);
assign l_7[9]    = ( l_8 [14] & !i[1707]) | ( l_8 [15] &  i[1707]);
assign l_7[10]    = (!l_8 [6] & !i[1707]) | ( l_8 [16] &  i[1707]);
assign l_7[11]    = ( l_8 [17] & !i[1707]) | ( l_8 [18] &  i[1707]);
assign l_7[12]    = (!l_8 [6] & !i[1707]) | (      i[1707]);
assign l_7[13]    = (!l_8 [9] & !i[1707]) | ( l_8 [19] &  i[1707]);
assign l_8[0]    = ( l_9 [0] & !i[1724]);
assign l_8[1]    = ( l_9 [1] & !i[1724]);
assign l_8[2]    = ( l_9 [2] & !i[1724]);
assign l_8[3]    = ( l_9 [3] & !i[1724]);
assign l_8[4]    = ( l_9 [4] & !i[1724]);
assign l_8[5]    = ( l_9 [5] & !i[1724]);
assign l_8[6]    = ( l_9 [6] & !i[1724]);
assign l_8[7]    = ( l_9 [7] & !i[1724]);
assign l_8[8]    = ( l_9 [8] & !i[1724]);
assign l_8[9]    = ( l_9 [9] & !i[1724]);
assign l_8[10]    = ( l_9 [10] & !i[1724]) | (      i[1724]);
assign l_8[11]    = ( l_9 [11] & !i[1724]) | (      i[1724]);
assign l_8[12]    = ( l_9 [12] & !i[1724]) | (      i[1724]);
assign l_8[13]    = ( l_9 [13] & !i[1724]) | (      i[1724]);
assign l_8[14]    = ( l_9 [14] & !i[1724]) | (      i[1724]);
assign l_8[15]    = ( l_9 [15] & !i[1724]) | (      i[1724]);
assign l_8[16]    = (!l_9 [5] & !i[1724]) | (      i[1724]);
assign l_8[17]    = ( l_9 [16] & !i[1724]) | (      i[1724]);
assign l_8[18]    = ( l_9 [17] & !i[1724]) | (      i[1724]);
assign l_8[19]    = (!l_9 [6] & !i[1724]) | (      i[1724]);
assign l_9[0]    = ( l_10 [0] & !i[1721]);
assign l_9[1]    = ( l_10 [1] & !i[1721]);
assign l_9[2]    = ( l_10 [2] & !i[1721]);
assign l_9[3]    = ( l_10 [3] & !i[1721]);
assign l_9[4]    = ( l_10 [4] & !i[1721]);
assign l_9[5]    = ( l_10 [5] & !i[1721]);
assign l_9[6]    = ( l_10 [6] & !i[1721]);
assign l_9[7]    = ( l_10 [7] & !i[1721]);
assign l_9[8]    = ( l_10 [8] & !i[1721]);
assign l_9[9]    = ( l_10 [9] & !i[1721]);
assign l_9[10]    = ( l_10 [10] & !i[1721]) | (      i[1721]);
assign l_9[11]    = ( l_10 [11] & !i[1721]) | (      i[1721]);
assign l_9[12]    = ( l_10 [12] & !i[1721]) | (      i[1721]);
assign l_9[13]    = ( l_10 [13] & !i[1721]) | (      i[1721]);
assign l_9[14]    = ( l_10 [14] & !i[1721]) | (      i[1721]);
assign l_9[15]    = ( l_10 [15] & !i[1721]) | (      i[1721]);
assign l_9[16]    = ( l_10 [16] & !i[1721]) | (      i[1721]);
assign l_9[17]    = ( l_10 [17] & !i[1721]) | (      i[1721]);
assign l_10[0]    = ( l_11 [0] &  i[1726]);
assign l_10[1]    = ( l_11 [1] &  i[1726]);
assign l_10[2]    = ( l_11 [2] &  i[1726]);
assign l_10[3]    = ( l_11 [3] &  i[1726]);
assign l_10[4]    = ( l_11 [4] &  i[1726]);
assign l_10[5]    = ( l_11 [5] &  i[1726]);
assign l_10[6]    = ( l_11 [6] &  i[1726]);
assign l_10[7]    = ( l_11 [7] &  i[1726]);
assign l_10[8]    = ( l_11 [8] &  i[1726]);
assign l_10[9]    = ( l_11 [9] &  i[1726]);
assign l_10[10]    = (!i[1726]) | ( l_11 [10] &  i[1726]);
assign l_10[11]    = (!i[1726]) | ( l_11 [11] &  i[1726]);
assign l_10[12]    = (!i[1726]) | ( l_11 [12] &  i[1726]);
assign l_10[13]    = (!i[1726]) | ( l_11 [13] &  i[1726]);
assign l_10[14]    = (!i[1726]) | ( l_11 [14] &  i[1726]);
assign l_10[15]    = (!i[1726]) | ( l_11 [15] &  i[1726]);
assign l_10[16]    = (!i[1726]) | ( l_11 [16] &  i[1726]);
assign l_10[17]    = (!i[1726]) | ( l_11 [17] &  i[1726]);
assign l_11[0]    = ( l_12 [0] &  i[1727]);
assign l_11[1]    = ( l_12 [1] &  i[1727]);
assign l_11[2]    = ( l_12 [2] &  i[1727]);
assign l_11[3]    = ( l_12 [3] &  i[1727]);
assign l_11[4]    = ( l_12 [4] &  i[1727]);
assign l_11[5]    = ( l_12 [5] &  i[1727]);
assign l_11[6]    = ( l_12 [6] &  i[1727]);
assign l_11[7]    = ( l_12 [7] &  i[1727]);
assign l_11[8]    = ( l_12 [8] &  i[1727]);
assign l_11[9]    = ( l_12 [9] &  i[1727]);
assign l_11[10]    = (!i[1727]) | ( l_12 [10] &  i[1727]);
assign l_11[11]    = (!i[1727]) | ( l_12 [11] &  i[1727]);
assign l_11[12]    = (!i[1727]) | ( l_12 [12] &  i[1727]);
assign l_11[13]    = (!i[1727]) | ( l_12 [13] &  i[1727]);
assign l_11[14]    = (!i[1727]) | ( l_12 [14] &  i[1727]);
assign l_11[15]    = (!i[1727]) | ( l_12 [15] &  i[1727]);
assign l_11[16]    = (!i[1727]) | ( l_12 [16] &  i[1727]);
assign l_11[17]    = (!i[1727]) | ( l_12 [17] &  i[1727]);
assign l_12[0]    = ( l_13 [0] & !i[1725]);
assign l_12[1]    = ( l_13 [1] & !i[1725]);
assign l_12[2]    = ( l_13 [2] & !i[1725]);
assign l_12[3]    = ( l_13 [3] & !i[1725]);
assign l_12[4]    = ( l_13 [4] & !i[1725]);
assign l_12[5]    = ( l_13 [5] & !i[1725]);
assign l_12[6]    = ( l_13 [6] & !i[1725]);
assign l_12[7]    = ( l_13 [7] & !i[1725]);
assign l_12[8]    = ( l_13 [8] & !i[1725]);
assign l_12[9]    = ( l_13 [9] & !i[1725]);
assign l_12[10]    = ( l_13 [10] & !i[1725]) | (      i[1725]);
assign l_12[11]    = ( l_13 [11] & !i[1725]) | (      i[1725]);
assign l_12[12]    = ( l_13 [12] & !i[1725]) | (      i[1725]);
assign l_12[13]    = ( l_13 [13] & !i[1725]) | (      i[1725]);
assign l_12[14]    = ( l_13 [14] & !i[1725]) | (      i[1725]);
assign l_12[15]    = ( l_13 [15] & !i[1725]) | (      i[1725]);
assign l_12[16]    = ( l_13 [16] & !i[1725]) | (      i[1725]);
assign l_12[17]    = ( l_13 [17] & !i[1725]) | (      i[1725]);
assign l_13[0]    = ( l_14 [0] & !i[1722]);
assign l_13[1]    = ( l_14 [1] & !i[1722]);
assign l_13[2]    = ( l_14 [2] & !i[1722]);
assign l_13[3]    = ( l_14 [3] & !i[1722]);
assign l_13[4]    = ( l_14 [4] & !i[1722]);
assign l_13[5]    = ( l_14 [5] & !i[1722]);
assign l_13[6]    = ( l_14 [6] & !i[1722]);
assign l_13[7]    = ( l_14 [7] & !i[1722]);
assign l_13[8]    = ( l_14 [8] & !i[1722]);
assign l_13[9]    = ( l_14 [9] & !i[1722]);
assign l_13[10]    = ( l_14 [10] & !i[1722]) | (      i[1722]);
assign l_13[11]    = ( l_14 [11] & !i[1722]) | (      i[1722]);
assign l_13[12]    = ( l_14 [12] & !i[1722]) | (      i[1722]);
assign l_13[13]    = ( l_14 [13] & !i[1722]) | (      i[1722]);
assign l_13[14]    = ( l_14 [14] & !i[1722]) | (      i[1722]);
assign l_13[15]    = ( l_14 [15] & !i[1722]) | (      i[1722]);
assign l_13[16]    = ( l_14 [16] & !i[1722]) | (      i[1722]);
assign l_13[17]    = ( l_14 [17] & !i[1722]) | (      i[1722]);
assign l_14[0]    = ( l_15 [0] & !i[1718]);
assign l_14[1]    = ( l_15 [1] & !i[1718]);
assign l_14[2]    = ( l_15 [2] & !i[1718]);
assign l_14[3]    = ( l_15 [3] & !i[1718]);
assign l_14[4]    = ( l_15 [4] & !i[1718]);
assign l_14[5]    = ( l_15 [5] & !i[1718]);
assign l_14[6]    = ( l_15 [6] & !i[1718]);
assign l_14[7]    = ( l_15 [7] & !i[1718]);
assign l_14[8]    = ( l_15 [8] & !i[1718]);
assign l_14[9]    = ( l_15 [9] & !i[1718]);
assign l_14[10]    = ( l_15 [10] & !i[1718]) | (      i[1718]);
assign l_14[11]    = ( l_15 [11] & !i[1718]) | (      i[1718]);
assign l_14[12]    = ( l_15 [12] & !i[1718]) | (      i[1718]);
assign l_14[13]    = ( l_15 [13] & !i[1718]) | (      i[1718]);
assign l_14[14]    = ( l_15 [14] & !i[1718]) | (      i[1718]);
assign l_14[15]    = ( l_15 [15] & !i[1718]) | (      i[1718]);
assign l_14[16]    = ( l_15 [16] & !i[1718]) | (      i[1718]);
assign l_14[17]    = ( l_15 [17] & !i[1718]) | (      i[1718]);
assign l_15[0]    = ( l_16 [0] & !i[1719]);
assign l_15[1]    = ( l_16 [1] & !i[1719]);
assign l_15[2]    = ( l_16 [2] & !i[1719]);
assign l_15[3]    = ( l_16 [3] & !i[1719]);
assign l_15[4]    = ( l_16 [4] & !i[1719]);
assign l_15[5]    = ( l_16 [5] & !i[1719]);
assign l_15[6]    = ( l_16 [6] & !i[1719]);
assign l_15[7]    = ( l_16 [7] & !i[1719]);
assign l_15[8]    = ( l_16 [8] & !i[1719]);
assign l_15[9]    = ( l_16 [9] & !i[1719]);
assign l_15[10]    = ( l_16 [10] & !i[1719]) | (      i[1719]);
assign l_15[11]    = ( l_16 [11] & !i[1719]) | (      i[1719]);
assign l_15[12]    = ( l_16 [12] & !i[1719]) | (      i[1719]);
assign l_15[13]    = ( l_16 [13] & !i[1719]) | (      i[1719]);
assign l_15[14]    = ( l_16 [14] & !i[1719]) | (      i[1719]);
assign l_15[15]    = ( l_16 [15] & !i[1719]) | (      i[1719]);
assign l_15[16]    = ( l_16 [16] & !i[1719]) | (      i[1719]);
assign l_15[17]    = ( l_16 [17] & !i[1719]) | (      i[1719]);
assign l_16[0]    = ( l_17 [0] &  i[1720]);
assign l_16[1]    = ( l_17 [1] &  i[1720]);
assign l_16[2]    = ( l_17 [2] &  i[1720]);
assign l_16[3]    = ( l_17 [3] &  i[1720]);
assign l_16[4]    = ( l_17 [4] &  i[1720]);
assign l_16[5]    = ( l_17 [5] &  i[1720]);
assign l_16[6]    = ( l_17 [6] &  i[1720]);
assign l_16[7]    = ( l_17 [7] &  i[1720]);
assign l_16[8]    = ( l_17 [8] &  i[1720]);
assign l_16[9]    =  i[1720];
assign l_16[10]    = (!i[1720]) | ( l_17 [9] &  i[1720]);
assign l_16[11]    = (!i[1720]) | ( l_17 [10] &  i[1720]);
assign l_16[12]    = (!i[1720]) | ( l_17 [1] &  i[1720]);
assign l_16[13]    = (!i[1720]) | ( l_17 [2] &  i[1720]);
assign l_16[14]    = (!i[1720]) | ( l_17 [3] &  i[1720]);
assign l_16[15]    = (!i[1720]) | ( l_17 [4] &  i[1720]);
assign l_16[16]    = (!i[1720]) | ( l_17 [11] &  i[1720]);
assign l_16[17]    = (!i[1720]) | ( l_17 [12] &  i[1720]);
assign l_17[0]    = ( l_18 [0] &  i[1829]);
assign l_17[1]    = ( l_18 [1]);
assign l_17[2]    = ( l_18 [2] & !i[1829]) | ( l_18 [1] &  i[1829]);
assign l_17[3]    = ( l_18 [3]);
assign l_17[4]    = ( l_18 [4] & !i[1829]) | ( l_18 [3] &  i[1829]);
assign l_17[5]    =  i[1829];
assign l_17[6]    = !i[1829];
assign l_17[7]    = ( l_18 [5] & !i[1829]) | ( l_18 [6] &  i[1829]);
assign l_17[8]    = ( l_18 [7]);
assign l_17[9]    = ( l_18 [8] & !i[1829]) | ( l_18 [9] &  i[1829]);
assign l_17[10]    = ( l_18 [8]);
assign l_17[11]    = ( l_18 [10] & !i[1829]) | ( l_18 [11] &  i[1829]);
assign l_17[12]    = ( l_18 [12]);
assign l_18[0]    = ( l_19 [0]);
assign l_18[1]    = ( l_19 [1] & !i[1798]) | ( l_19 [2] &  i[1798]);
assign l_18[2]    = ( l_19 [3] & !i[1798]) | ( l_19 [4] &  i[1798]);
assign l_18[3]    = ( l_19 [5] & !i[1798]) | ( l_19 [6] &  i[1798]);
assign l_18[4]    = ( l_19 [7] & !i[1798]) | ( l_19 [8] &  i[1798]);
assign l_18[5]    = ( l_19 [9]);
assign l_18[6]    = ( l_19 [10]);
assign l_18[7]    = ( l_19 [11] & !i[1798]) | ( l_19 [12] &  i[1798]);
assign l_18[8]    = ( l_19 [13]);
assign l_18[9]    = ( l_19 [14]);
assign l_18[10]    = ( l_19 [15]);
assign l_18[11]    = ( l_19 [16]);
assign l_18[12]    = ( l_19 [17] & !i[1798]) | ( l_19 [18] &  i[1798]);
assign l_19[0]    = ( l_20 [0]);
assign l_19[1]    = ( l_20 [1] & !i[1809]);
assign l_19[2]    = (!i[1809]) | ( l_20 [2] &  i[1809]);
assign l_19[3]    = ( l_20 [3] & !i[1809]);
assign l_19[4]    = (!i[1809]) | ( l_20 [4] &  i[1809]);
assign l_19[5]    = ( l_20 [5] & !i[1809]) | ( l_20 [6] &  i[1809]);
assign l_19[6]    = ( l_20 [6] & !i[1809]) | ( l_20 [7] &  i[1809]);
assign l_19[7]    = ( l_20 [8] & !i[1809]) | ( l_20 [6] &  i[1809]);
assign l_19[8]    = ( l_20 [6] & !i[1809]) | ( l_20 [9] &  i[1809]);
assign l_19[9]    = ( l_20 [10] & !i[1809]) | ( l_20 [11] &  i[1809]);
assign l_19[10]    = ( l_20 [12] & !i[1809]) | ( l_20 [13] &  i[1809]);
assign l_19[11]    = ( l_20 [14]);
assign l_19[12]    = ( l_20 [15]);
assign l_19[13]    = ( l_20 [16]);
assign l_19[14]    = ( l_20 [17]);
assign l_19[15]    = ( l_20 [18] & !i[1809]) | ( l_20 [19] &  i[1809]);
assign l_19[16]    = ( l_20 [20] & !i[1809]) | ( l_20 [21] &  i[1809]);
assign l_19[17]    = ( l_20 [22]);
assign l_19[18]    = ( l_20 [23]);

endmodule
