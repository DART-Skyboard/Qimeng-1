module module_output_bit_63(i,o);

input [1893:0] i;
output  o;

wire [0:0] l_0;
wire [1:0] l_1;
wire [3:0] l_2;
wire [7:0] l_3;
wire [13:0] l_4;
wire [13:0] l_5;
wire [13:0] l_6;
wire [13:0] l_7;
wire [19:0] l_8;
wire [17:0] l_9;
wire [17:0] l_10;
wire [17:0] l_11;
wire [17:0] l_12;
wire [17:0] l_13;
wire [17:0] l_14;
wire [17:0] l_15;
wire [17:0] l_16;
wire [12:0] l_17;
wire [12:0] l_18;
wire [18:0] l_19;
wire [23:0] l_20;
wire [23:0] l_21;
wire [27:0] l_22;
wire [35:0] l_23;
wire [51:0] l_24;
wire [53:0] l_25;
wire [85:0] l_26;
wire [89:0] l_27;
wire [97:0] l_28;
wire [113:0] l_29;
wire [145:0] l_30;

assign	l_30[145:0]	= 146'b0;

assign o = l_0[0];

assign l_0[0]    = ( l_1 [0] & !i[63]) | ( l_1 [1] &  i[63]);
assign l_1[0]    = ( l_2 [0] & !i[1713]) | ( l_2 [1] &  i[1713]);
assign l_1[1]    = ( l_2 [2] & !i[1713]) | ( l_2 [3] &  i[1713]);
assign l_2[0]    = ( l_3 [0] & !i[1714]) | ( l_3 [1] &  i[1714]);
assign l_2[1]    = ( l_3 [2] & !i[1714]) | ( l_3 [3] &  i[1714]);
assign l_2[2]    = ( l_3 [4] & !i[1714]) | ( l_3 [5] &  i[1714]);
assign l_2[3]    = ( l_3 [6] & !i[1714]) | ( l_3 [7] &  i[1714]);
assign l_3[0]    = ( l_4 [0] &  i[1715]);
assign l_3[1]    = ( l_4 [1] & !i[1715]) | ( l_4 [2] &  i[1715]);
assign l_3[2]    = ( l_4 [3] & !i[1715]) | ( l_4 [4] &  i[1715]);
assign l_3[3]    = ( l_4 [5] & !i[1715]) | ( l_4 [6] &  i[1715]);
assign l_3[4]    = (!i[1715]) | ( l_4 [7] &  i[1715]);
assign l_3[5]    = ( l_4 [8] & !i[1715]) | ( l_4 [9] &  i[1715]);
assign l_3[6]    = ( l_4 [10] & !i[1715]) | ( l_4 [11] &  i[1715]);
assign l_3[7]    = ( l_4 [12] & !i[1715]) | ( l_4 [13] &  i[1715]);
assign l_4[0]    = ( l_5 [0] & !i[1716]);
assign l_4[1]    = ( l_5 [1] & !i[1716]);
assign l_4[2]    = ( l_5 [2] & !i[1716]);
assign l_4[3]    = ( l_5 [3] & !i[1716]);
assign l_4[4]    = ( l_5 [4] & !i[1716]);
assign l_4[5]    = ( l_5 [5] & !i[1716]);
assign l_4[6]    = ( l_5 [6] & !i[1716]);
assign l_4[7]    = ( l_5 [7] & !i[1716]) | (      i[1716]);
assign l_4[8]    = ( l_5 [8] & !i[1716]) | (      i[1716]);
assign l_4[9]    = ( l_5 [9] & !i[1716]) | (      i[1716]);
assign l_4[10]    = ( l_5 [10] & !i[1716]) | (      i[1716]);
assign l_4[11]    = ( l_5 [11] & !i[1716]) | (      i[1716]);
assign l_4[12]    = ( l_5 [12] & !i[1716]) | (      i[1716]);
assign l_4[13]    = ( l_5 [13] & !i[1716]) | (      i[1716]);
assign l_5[0]    = ( l_6 [0] & !i[1717]);
assign l_5[1]    = ( l_6 [1] & !i[1717]);
assign l_5[2]    = ( l_6 [2] & !i[1717]);
assign l_5[3]    = ( l_6 [3] & !i[1717]);
assign l_5[4]    = ( l_6 [4] & !i[1717]);
assign l_5[5]    = ( l_6 [5] & !i[1717]);
assign l_5[6]    = ( l_6 [6] & !i[1717]);
assign l_5[7]    = ( l_6 [7] & !i[1717]) | (      i[1717]);
assign l_5[8]    = ( l_6 [8] & !i[1717]) | (      i[1717]);
assign l_5[9]    = ( l_6 [9] & !i[1717]) | (      i[1717]);
assign l_5[10]    = ( l_6 [10] & !i[1717]) | (      i[1717]);
assign l_5[11]    = ( l_6 [11] & !i[1717]) | (      i[1717]);
assign l_5[12]    = ( l_6 [12] & !i[1717]) | (      i[1717]);
assign l_5[13]    = ( l_6 [13] & !i[1717]) | (      i[1717]);
assign l_6[0]    = ( l_7 [0] &  i[1723]);
assign l_6[1]    = ( l_7 [1] &  i[1723]);
assign l_6[2]    = ( l_7 [2] &  i[1723]);
assign l_6[3]    = ( l_7 [3] &  i[1723]);
assign l_6[4]    = ( l_7 [4] &  i[1723]);
assign l_6[5]    = ( l_7 [5] &  i[1723]);
assign l_6[6]    = ( l_7 [6] &  i[1723]);
assign l_6[7]    = (!i[1723]) | ( l_7 [7] &  i[1723]);
assign l_6[8]    = (!i[1723]) | ( l_7 [8] &  i[1723]);
assign l_6[9]    = (!i[1723]) | ( l_7 [9] &  i[1723]);
assign l_6[10]    = (!i[1723]) | ( l_7 [10] &  i[1723]);
assign l_6[11]    = (!i[1723]) | ( l_7 [11] &  i[1723]);
assign l_6[12]    = (!i[1723]) | ( l_7 [12] &  i[1723]);
assign l_6[13]    = (!i[1723]) | ( l_7 [13] &  i[1723]);
assign l_7[0]    = ( l_8 [0] & !i[1707]);
assign l_7[1]    = ( l_8 [1] & !i[1707]) | ( l_8 [2] &  i[1707]);
assign l_7[2]    = ( l_8 [3] & !i[1707]) | ( l_8 [4] &  i[1707]);
assign l_7[3]    = ( l_8 [5] & !i[1707]) | ( l_8 [6] &  i[1707]);
assign l_7[4]    = ( l_8 [7] & !i[1707]) | ( l_8 [8] &  i[1707]);
assign l_7[5]    = ( l_8 [5] & !i[1707]) | ( l_8 [9] &  i[1707]);
assign l_7[6]    = ( l_8 [5] &  i[1707]);
assign l_7[7]    = ( l_8 [10] & !i[1707]) | ( l_8 [11] &  i[1707]);
assign l_7[8]    = ( l_8 [12] & !i[1707]) | ( l_8 [13] &  i[1707]);
assign l_7[9]    = ( l_8 [14] & !i[1707]) | ( l_8 [15] &  i[1707]);
assign l_7[10]    = (!l_8 [6] & !i[1707]) | ( l_8 [16] &  i[1707]);
assign l_7[11]    = ( l_8 [17] & !i[1707]) | ( l_8 [18] &  i[1707]);
assign l_7[12]    = (!l_8 [6] & !i[1707]) | (      i[1707]);
assign l_7[13]    = (!l_8 [9] & !i[1707]) | ( l_8 [19] &  i[1707]);
assign l_8[0]    = ( l_9 [0] & !i[1724]);
assign l_8[1]    = ( l_9 [1] & !i[1724]);
assign l_8[2]    = ( l_9 [2] & !i[1724]);
assign l_8[3]    = ( l_9 [3] & !i[1724]);
assign l_8[4]    = ( l_9 [4] & !i[1724]);
assign l_8[5]    = ( l_9 [5] & !i[1724]);
assign l_8[6]    = ( l_9 [6] & !i[1724]);
assign l_8[7]    = ( l_9 [7] & !i[1724]);
assign l_8[8]    = ( l_9 [8] & !i[1724]);
assign l_8[9]    = ( l_9 [9] & !i[1724]);
assign l_8[10]    = ( l_9 [10] & !i[1724]) | (      i[1724]);
assign l_8[11]    = ( l_9 [11] & !i[1724]) | (      i[1724]);
assign l_8[12]    = ( l_9 [12] & !i[1724]) | (      i[1724]);
assign l_8[13]    = ( l_9 [13] & !i[1724]) | (      i[1724]);
assign l_8[14]    = ( l_9 [14] & !i[1724]) | (      i[1724]);
assign l_8[15]    = ( l_9 [15] & !i[1724]) | (      i[1724]);
assign l_8[16]    = (!l_9 [5] & !i[1724]) | (      i[1724]);
assign l_8[17]    = ( l_9 [16] & !i[1724]) | (      i[1724]);
assign l_8[18]    = ( l_9 [17] & !i[1724]) | (      i[1724]);
assign l_8[19]    = (!l_9 [6] & !i[1724]) | (      i[1724]);
assign l_9[0]    = ( l_10 [0] & !i[1721]);
assign l_9[1]    = ( l_10 [1] & !i[1721]);
assign l_9[2]    = ( l_10 [2] & !i[1721]);
assign l_9[3]    = ( l_10 [3] & !i[1721]);
assign l_9[4]    = ( l_10 [4] & !i[1721]);
assign l_9[5]    = ( l_10 [5] & !i[1721]);
assign l_9[6]    = ( l_10 [6] & !i[1721]);
assign l_9[7]    = ( l_10 [7] & !i[1721]);
assign l_9[8]    = ( l_10 [8] & !i[1721]);
assign l_9[9]    = ( l_10 [9] & !i[1721]);
assign l_9[10]    = ( l_10 [10] & !i[1721]) | (      i[1721]);
assign l_9[11]    = ( l_10 [11] & !i[1721]) | (      i[1721]);
assign l_9[12]    = ( l_10 [12] & !i[1721]) | (      i[1721]);
assign l_9[13]    = ( l_10 [13] & !i[1721]) | (      i[1721]);
assign l_9[14]    = ( l_10 [14] & !i[1721]) | (      i[1721]);
assign l_9[15]    = ( l_10 [15] & !i[1721]) | (      i[1721]);
assign l_9[16]    = ( l_10 [16] & !i[1721]) | (      i[1721]);
assign l_9[17]    = ( l_10 [17] & !i[1721]) | (      i[1721]);
assign l_10[0]    = ( l_11 [0] &  i[1726]);
assign l_10[1]    = ( l_11 [1] &  i[1726]);
assign l_10[2]    = ( l_11 [2] &  i[1726]);
assign l_10[3]    = ( l_11 [3] &  i[1726]);
assign l_10[4]    = ( l_11 [4] &  i[1726]);
assign l_10[5]    = ( l_11 [5] &  i[1726]);
assign l_10[6]    = ( l_11 [6] &  i[1726]);
assign l_10[7]    = ( l_11 [7] &  i[1726]);
assign l_10[8]    = ( l_11 [8] &  i[1726]);
assign l_10[9]    = ( l_11 [9] &  i[1726]);
assign l_10[10]    = (!i[1726]) | ( l_11 [10] &  i[1726]);
assign l_10[11]    = (!i[1726]) | ( l_11 [11] &  i[1726]);
assign l_10[12]    = (!i[1726]) | ( l_11 [12] &  i[1726]);
assign l_10[13]    = (!i[1726]) | ( l_11 [13] &  i[1726]);
assign l_10[14]    = (!i[1726]) | ( l_11 [14] &  i[1726]);
assign l_10[15]    = (!i[1726]) | ( l_11 [15] &  i[1726]);
assign l_10[16]    = (!i[1726]) | ( l_11 [16] &  i[1726]);
assign l_10[17]    = (!i[1726]) | ( l_11 [17] &  i[1726]);
assign l_11[0]    = ( l_12 [0] &  i[1727]);
assign l_11[1]    = ( l_12 [1] &  i[1727]);
assign l_11[2]    = ( l_12 [2] &  i[1727]);
assign l_11[3]    = ( l_12 [3] &  i[1727]);
assign l_11[4]    = ( l_12 [4] &  i[1727]);
assign l_11[5]    = ( l_12 [5] &  i[1727]);
assign l_11[6]    = ( l_12 [6] &  i[1727]);
assign l_11[7]    = ( l_12 [7] &  i[1727]);
assign l_11[8]    = ( l_12 [8] &  i[1727]);
assign l_11[9]    = ( l_12 [9] &  i[1727]);
assign l_11[10]    = (!i[1727]) | ( l_12 [10] &  i[1727]);
assign l_11[11]    = (!i[1727]) | ( l_12 [11] &  i[1727]);
assign l_11[12]    = (!i[1727]) | ( l_12 [12] &  i[1727]);
assign l_11[13]    = (!i[1727]) | ( l_12 [13] &  i[1727]);
assign l_11[14]    = (!i[1727]) | ( l_12 [14] &  i[1727]);
assign l_11[15]    = (!i[1727]) | ( l_12 [15] &  i[1727]);
assign l_11[16]    = (!i[1727]) | ( l_12 [16] &  i[1727]);
assign l_11[17]    = (!i[1727]) | ( l_12 [17] &  i[1727]);
assign l_12[0]    = ( l_13 [0] & !i[1725]);
assign l_12[1]    = ( l_13 [1] & !i[1725]);
assign l_12[2]    = ( l_13 [2] & !i[1725]);
assign l_12[3]    = ( l_13 [3] & !i[1725]);
assign l_12[4]    = ( l_13 [4] & !i[1725]);
assign l_12[5]    = ( l_13 [5] & !i[1725]);
assign l_12[6]    = ( l_13 [6] & !i[1725]);
assign l_12[7]    = ( l_13 [7] & !i[1725]);
assign l_12[8]    = ( l_13 [8] & !i[1725]);
assign l_12[9]    = ( l_13 [9] & !i[1725]);
assign l_12[10]    = ( l_13 [10] & !i[1725]) | (      i[1725]);
assign l_12[11]    = ( l_13 [11] & !i[1725]) | (      i[1725]);
assign l_12[12]    = ( l_13 [12] & !i[1725]) | (      i[1725]);
assign l_12[13]    = ( l_13 [13] & !i[1725]) | (      i[1725]);
assign l_12[14]    = ( l_13 [14] & !i[1725]) | (      i[1725]);
assign l_12[15]    = ( l_13 [15] & !i[1725]) | (      i[1725]);
assign l_12[16]    = ( l_13 [16] & !i[1725]) | (      i[1725]);
assign l_12[17]    = ( l_13 [17] & !i[1725]) | (      i[1725]);
assign l_13[0]    = ( l_14 [0] & !i[1722]);
assign l_13[1]    = ( l_14 [1] & !i[1722]);
assign l_13[2]    = ( l_14 [2] & !i[1722]);
assign l_13[3]    = ( l_14 [3] & !i[1722]);
assign l_13[4]    = ( l_14 [4] & !i[1722]);
assign l_13[5]    = ( l_14 [5] & !i[1722]);
assign l_13[6]    = ( l_14 [6] & !i[1722]);
assign l_13[7]    = ( l_14 [7] & !i[1722]);
assign l_13[8]    = ( l_14 [8] & !i[1722]);
assign l_13[9]    = ( l_14 [9] & !i[1722]);
assign l_13[10]    = ( l_14 [10] & !i[1722]) | (      i[1722]);
assign l_13[11]    = ( l_14 [11] & !i[1722]) | (      i[1722]);
assign l_13[12]    = ( l_14 [12] & !i[1722]) | (      i[1722]);
assign l_13[13]    = ( l_14 [13] & !i[1722]) | (      i[1722]);
assign l_13[14]    = ( l_14 [14] & !i[1722]) | (      i[1722]);
assign l_13[15]    = ( l_14 [15] & !i[1722]) | (      i[1722]);
assign l_13[16]    = ( l_14 [16] & !i[1722]) | (      i[1722]);
assign l_13[17]    = ( l_14 [17] & !i[1722]) | (      i[1722]);
assign l_14[0]    = ( l_15 [0] & !i[1718]);
assign l_14[1]    = ( l_15 [1] & !i[1718]);
assign l_14[2]    = ( l_15 [2] & !i[1718]);
assign l_14[3]    = ( l_15 [3] & !i[1718]);
assign l_14[4]    = ( l_15 [4] & !i[1718]);
assign l_14[5]    = ( l_15 [5] & !i[1718]);
assign l_14[6]    = ( l_15 [6] & !i[1718]);
assign l_14[7]    = ( l_15 [7] & !i[1718]);
assign l_14[8]    = ( l_15 [8] & !i[1718]);
assign l_14[9]    = ( l_15 [9] & !i[1718]);
assign l_14[10]    = ( l_15 [10] & !i[1718]) | (      i[1718]);
assign l_14[11]    = ( l_15 [11] & !i[1718]) | (      i[1718]);
assign l_14[12]    = ( l_15 [12] & !i[1718]) | (      i[1718]);
assign l_14[13]    = ( l_15 [13] & !i[1718]) | (      i[1718]);
assign l_14[14]    = ( l_15 [14] & !i[1718]) | (      i[1718]);
assign l_14[15]    = ( l_15 [15] & !i[1718]) | (      i[1718]);
assign l_14[16]    = ( l_15 [16] & !i[1718]) | (      i[1718]);
assign l_14[17]    = ( l_15 [17] & !i[1718]) | (      i[1718]);
assign l_15[0]    = ( l_16 [0] & !i[1719]);
assign l_15[1]    = ( l_16 [1] & !i[1719]);
assign l_15[2]    = ( l_16 [2] & !i[1719]);
assign l_15[3]    = ( l_16 [3] & !i[1719]);
assign l_15[4]    = ( l_16 [4] & !i[1719]);
assign l_15[5]    = ( l_16 [5] & !i[1719]);
assign l_15[6]    = ( l_16 [6] & !i[1719]);
assign l_15[7]    = ( l_16 [7] & !i[1719]);
assign l_15[8]    = ( l_16 [8] & !i[1719]);
assign l_15[9]    = ( l_16 [9] & !i[1719]);
assign l_15[10]    = ( l_16 [10] & !i[1719]) | (      i[1719]);
assign l_15[11]    = ( l_16 [11] & !i[1719]) | (      i[1719]);
assign l_15[12]    = ( l_16 [12] & !i[1719]) | (      i[1719]);
assign l_15[13]    = ( l_16 [13] & !i[1719]) | (      i[1719]);
assign l_15[14]    = ( l_16 [14] & !i[1719]) | (      i[1719]);
assign l_15[15]    = ( l_16 [15] & !i[1719]) | (      i[1719]);
assign l_15[16]    = ( l_16 [16] & !i[1719]) | (      i[1719]);
assign l_15[17]    = ( l_16 [17] & !i[1719]) | (      i[1719]);
assign l_16[0]    = ( l_17 [0] &  i[1720]);
assign l_16[1]    = ( l_17 [1] &  i[1720]);
assign l_16[2]    = ( l_17 [2] &  i[1720]);
assign l_16[3]    = ( l_17 [3] &  i[1720]);
assign l_16[4]    = ( l_17 [4] &  i[1720]);
assign l_16[5]    = ( l_17 [5] &  i[1720]);
assign l_16[6]    = ( l_17 [6] &  i[1720]);
assign l_16[7]    = ( l_17 [7] &  i[1720]);
assign l_16[8]    = ( l_17 [8] &  i[1720]);
assign l_16[9]    =  i[1720];
assign l_16[10]    = (!i[1720]) | ( l_17 [9] &  i[1720]);
assign l_16[11]    = (!i[1720]) | ( l_17 [10] &  i[1720]);
assign l_16[12]    = (!i[1720]) | ( l_17 [1] &  i[1720]);
assign l_16[13]    = (!i[1720]) | ( l_17 [2] &  i[1720]);
assign l_16[14]    = (!i[1720]) | ( l_17 [3] &  i[1720]);
assign l_16[15]    = (!i[1720]) | ( l_17 [4] &  i[1720]);
assign l_16[16]    = (!i[1720]) | ( l_17 [11] &  i[1720]);
assign l_16[17]    = (!i[1720]) | ( l_17 [12] &  i[1720]);
assign l_17[0]    = ( l_18 [0] &  i[1829]);
assign l_17[1]    = ( l_18 [1]);
assign l_17[2]    = ( l_18 [2] & !i[1829]) | ( l_18 [1] &  i[1829]);
assign l_17[3]    = ( l_18 [3]);
assign l_17[4]    = ( l_18 [4] & !i[1829]) | ( l_18 [3] &  i[1829]);
assign l_17[5]    =  i[1829];
assign l_17[6]    = !i[1829];
assign l_17[7]    = ( l_18 [5] & !i[1829]) | ( l_18 [6] &  i[1829]);
assign l_17[8]    = ( l_18 [7]);
assign l_17[9]    = ( l_18 [8] & !i[1829]) | ( l_18 [9] &  i[1829]);
assign l_17[10]    = ( l_18 [8]);
assign l_17[11]    = ( l_18 [10] & !i[1829]) | ( l_18 [11] &  i[1829]);
assign l_17[12]    = ( l_18 [12]);
assign l_18[0]    = ( l_19 [0]);
assign l_18[1]    = ( l_19 [1] & !i[1798]) | ( l_19 [2] &  i[1798]);
assign l_18[2]    = ( l_19 [3] & !i[1798]) | ( l_19 [4] &  i[1798]);
assign l_18[3]    = ( l_19 [5] & !i[1798]) | ( l_19 [6] &  i[1798]);
assign l_18[4]    = ( l_19 [7] & !i[1798]) | ( l_19 [8] &  i[1798]);
assign l_18[5]    = ( l_19 [9]);
assign l_18[6]    = ( l_19 [10]);
assign l_18[7]    = ( l_19 [11] & !i[1798]) | ( l_19 [12] &  i[1798]);
assign l_18[8]    = ( l_19 [13]);
assign l_18[9]    = ( l_19 [14]);
assign l_18[10]    = ( l_19 [15]);
assign l_18[11]    = ( l_19 [16]);
assign l_18[12]    = ( l_19 [17] & !i[1798]) | ( l_19 [18] &  i[1798]);
assign l_19[0]    = ( l_20 [0]);
assign l_19[1]    = ( l_20 [1] & !i[1809]);
assign l_19[2]    = (!i[1809]) | ( l_20 [2] &  i[1809]);
assign l_19[3]    = ( l_20 [3] & !i[1809]);
assign l_19[4]    = (!i[1809]) | ( l_20 [4] &  i[1809]);
assign l_19[5]    = ( l_20 [5] & !i[1809]) | ( l_20 [6] &  i[1809]);
assign l_19[6]    = ( l_20 [6] & !i[1809]) | ( l_20 [7] &  i[1809]);
assign l_19[7]    = ( l_20 [8] & !i[1809]) | ( l_20 [6] &  i[1809]);
assign l_19[8]    = ( l_20 [6] & !i[1809]) | ( l_20 [9] &  i[1809]);
assign l_19[9]    = ( l_20 [10] & !i[1809]) | ( l_20 [11] &  i[1809]);
assign l_19[10]    = ( l_20 [12] & !i[1809]) | ( l_20 [13] &  i[1809]);
assign l_19[11]    = ( l_20 [14]);
assign l_19[12]    = ( l_20 [15]);
assign l_19[13]    = ( l_20 [16]);
assign l_19[14]    = ( l_20 [17]);
assign l_19[15]    = ( l_20 [18] & !i[1809]) | ( l_20 [19] &  i[1809]);
assign l_19[16]    = ( l_20 [20] & !i[1809]) | ( l_20 [21] &  i[1809]);
assign l_19[17]    = ( l_20 [22]);
assign l_19[18]    = ( l_20 [23]);
assign l_20[0]    = ( l_21 [0] & !i[1702]);
assign l_20[1]    = ( l_21 [1] & !i[1702]) | ( l_21 [2] &  i[1702]);
assign l_20[2]    = ( l_21 [3] & !i[1702]) | ( l_21 [4] &  i[1702]);
assign l_20[3]    = ( l_21 [5] & !i[1702]) | ( l_21 [6] &  i[1702]);
assign l_20[4]    = ( l_21 [7] & !i[1702]) | ( l_21 [8] &  i[1702]);
assign l_20[5]    = ( l_21 [9] & !i[1702]) | ( l_21 [10] &  i[1702]);
assign l_20[6]    = ( l_21 [11]);
assign l_20[7]    = ( l_21 [12] & !i[1702]) | ( l_21 [13] &  i[1702]);
assign l_20[8]    = ( l_21 [14] & !i[1702]) | ( l_21 [15] &  i[1702]);
assign l_20[9]    = ( l_21 [16] & !i[1702]) | ( l_21 [17] &  i[1702]);
assign l_20[10]    = ( l_21 [18] & !i[1702]);
assign l_20[11]    = ( l_21 [19] & !i[1702]);
assign l_20[12]    = ( l_21 [20] & !i[1702]);
assign l_20[13]    = ( l_21 [21] & !i[1702]);
assign l_20[14]    = ( l_21 [22] & !i[1702]);
assign l_20[15]    = ( l_21 [23] & !i[1702]);
assign l_20[16]    =  i[1702];
assign l_20[17]    = ( l_21 [0] & !i[1702]) | (      i[1702]);
assign l_20[18]    = ( l_21 [18] & !i[1702]) | (      i[1702]);
assign l_20[19]    = ( l_21 [19] & !i[1702]) | (      i[1702]);
assign l_20[20]    = ( l_21 [20] & !i[1702]) | (      i[1702]);
assign l_20[21]    = ( l_21 [21] & !i[1702]) | (      i[1702]);
assign l_20[22]    = ( l_21 [22] & !i[1702]) | (      i[1702]);
assign l_20[23]    = ( l_21 [23] & !i[1702]) | (      i[1702]);
assign l_21[0]    = ( l_22 [0]);
assign l_21[1]    = ( l_22 [1] & !i[1803]);
assign l_21[2]    = ( l_22 [2] & !i[1803]);
assign l_21[3]    = (!i[1803]) | ( l_22 [3] &  i[1803]);
assign l_21[4]    = (!i[1803]) | ( l_22 [4] &  i[1803]);
assign l_21[5]    = ( l_22 [5] & !i[1803]);
assign l_21[6]    = ( l_22 [6] & !i[1803]);
assign l_21[7]    = (!i[1803]) | ( l_22 [7] &  i[1803]);
assign l_21[8]    = (!i[1803]) | ( l_22 [8] &  i[1803]);
assign l_21[9]    = ( l_22 [9] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[10]    = ( l_22 [11] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[11]    = ( l_22 [10]);
assign l_21[12]    = ( l_22 [10] & !i[1803]) | ( l_22 [12] &  i[1803]);
assign l_21[13]    = ( l_22 [10] & !i[1803]) | ( l_22 [13] &  i[1803]);
assign l_21[14]    = ( l_22 [14] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[15]    = ( l_22 [15] & !i[1803]) | ( l_22 [10] &  i[1803]);
assign l_21[16]    = ( l_22 [10] & !i[1803]) | ( l_22 [16] &  i[1803]);
assign l_21[17]    = ( l_22 [10] & !i[1803]) | ( l_22 [17] &  i[1803]);
assign l_21[18]    = ( l_22 [18] & !i[1803]) | ( l_22 [19] &  i[1803]);
assign l_21[19]    = ( l_22 [20] & !i[1803]) | ( l_22 [21] &  i[1803]);
assign l_21[20]    = ( l_22 [22] & !i[1803]) | ( l_22 [23] &  i[1803]);
assign l_21[21]    = ( l_22 [24] & !i[1803]) | ( l_22 [25] &  i[1803]);
assign l_21[22]    = ( l_22 [26]);
assign l_21[23]    = ( l_22 [27]);
assign l_22[0]    = ( l_23 [0]);
assign l_22[1]    = ( l_23 [1] & !i[1801]);
assign l_22[2]    = ( l_23 [2] & !i[1801]);
assign l_22[3]    = (!i[1801]) | ( l_23 [3] &  i[1801]);
assign l_22[4]    = (!i[1801]) | ( l_23 [4] &  i[1801]);
assign l_22[5]    = ( l_23 [5] & !i[1801]);
assign l_22[6]    = ( l_23 [6] & !i[1801]);
assign l_22[7]    = (!i[1801]) | ( l_23 [7] &  i[1801]);
assign l_22[8]    = (!i[1801]) | ( l_23 [8] &  i[1801]);
assign l_22[9]    = ( l_23 [9] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[10]    = ( l_23 [10]);
assign l_22[11]    = ( l_23 [11] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[12]    = ( l_23 [10] & !i[1801]) | ( l_23 [12] &  i[1801]);
assign l_22[13]    = ( l_23 [10] & !i[1801]) | ( l_23 [13] &  i[1801]);
assign l_22[14]    = ( l_23 [14] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[15]    = ( l_23 [15] & !i[1801]) | ( l_23 [10] &  i[1801]);
assign l_22[16]    = ( l_23 [10] & !i[1801]) | ( l_23 [16] &  i[1801]);
assign l_22[17]    = ( l_23 [10] & !i[1801]) | ( l_23 [17] &  i[1801]);
assign l_22[18]    = ( l_23 [18] & !i[1801]) | ( l_23 [19] &  i[1801]);
assign l_22[19]    = ( l_23 [20] & !i[1801]) | ( l_23 [21] &  i[1801]);
assign l_22[20]    = ( l_23 [22] & !i[1801]) | ( l_23 [23] &  i[1801]);
assign l_22[21]    = ( l_23 [24] & !i[1801]) | ( l_23 [25] &  i[1801]);
assign l_22[22]    = ( l_23 [26] & !i[1801]) | ( l_23 [27] &  i[1801]);
assign l_22[23]    = ( l_23 [28] & !i[1801]) | ( l_23 [29] &  i[1801]);
assign l_22[24]    = ( l_23 [30] & !i[1801]) | ( l_23 [31] &  i[1801]);
assign l_22[25]    = ( l_23 [32] & !i[1801]) | ( l_23 [33] &  i[1801]);
assign l_22[26]    = ( l_23 [34]);
assign l_22[27]    = ( l_23 [35]);
assign l_23[0]    = ( l_24 [0]);
assign l_23[1]    = ( l_24 [1] & !i[1805]);
assign l_23[2]    = ( l_24 [2] & !i[1805]);
assign l_23[3]    = (!i[1805]) | ( l_24 [3] &  i[1805]);
assign l_23[4]    = (!i[1805]) | ( l_24 [4] &  i[1805]);
assign l_23[5]    = ( l_24 [5] & !i[1805]);
assign l_23[6]    = ( l_24 [6] & !i[1805]);
assign l_23[7]    = (!i[1805]) | ( l_24 [7] &  i[1805]);
assign l_23[8]    = (!i[1805]) | ( l_24 [8] &  i[1805]);
assign l_23[9]    = ( l_24 [9] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[10]    = ( l_24 [10]);
assign l_23[11]    = ( l_24 [11] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[12]    = ( l_24 [10] & !i[1805]) | ( l_24 [12] &  i[1805]);
assign l_23[13]    = ( l_24 [10] & !i[1805]) | ( l_24 [13] &  i[1805]);
assign l_23[14]    = ( l_24 [14] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[15]    = ( l_24 [15] & !i[1805]) | ( l_24 [10] &  i[1805]);
assign l_23[16]    = ( l_24 [10] & !i[1805]) | ( l_24 [16] &  i[1805]);
assign l_23[17]    = ( l_24 [10] & !i[1805]) | ( l_24 [17] &  i[1805]);
assign l_23[18]    = ( l_24 [18] & !i[1805]) | ( l_24 [19] &  i[1805]);
assign l_23[19]    = ( l_24 [20] & !i[1805]) | ( l_24 [21] &  i[1805]);
assign l_23[20]    = ( l_24 [22] & !i[1805]) | ( l_24 [23] &  i[1805]);
assign l_23[21]    = ( l_24 [24] & !i[1805]) | ( l_24 [25] &  i[1805]);
assign l_23[22]    = ( l_24 [26] & !i[1805]) | ( l_24 [27] &  i[1805]);
assign l_23[23]    = ( l_24 [28] & !i[1805]) | ( l_24 [29] &  i[1805]);
assign l_23[24]    = ( l_24 [30] & !i[1805]) | ( l_24 [31] &  i[1805]);
assign l_23[25]    = ( l_24 [32] & !i[1805]) | ( l_24 [33] &  i[1805]);
assign l_23[26]    = ( l_24 [34] & !i[1805]) | ( l_24 [35] &  i[1805]);
assign l_23[27]    = ( l_24 [36] & !i[1805]) | ( l_24 [37] &  i[1805]);
assign l_23[28]    = ( l_24 [38] & !i[1805]) | ( l_24 [39] &  i[1805]);
assign l_23[29]    = ( l_24 [40] & !i[1805]) | ( l_24 [41] &  i[1805]);
assign l_23[30]    = ( l_24 [42] & !i[1805]) | ( l_24 [43] &  i[1805]);
assign l_23[31]    = ( l_24 [44] & !i[1805]) | ( l_24 [45] &  i[1805]);
assign l_23[32]    = ( l_24 [46] & !i[1805]) | ( l_24 [47] &  i[1805]);
assign l_23[33]    = ( l_24 [48] & !i[1805]) | ( l_24 [49] &  i[1805]);
assign l_23[34]    = ( l_24 [50]);
assign l_23[35]    = ( l_24 [51]);
assign l_24[0]    = ( l_25 [0]);
assign l_24[1]    = ( l_25 [1] & !i[1808]);
assign l_24[2]    = ( l_25 [2] & !i[1808]);
assign l_24[3]    = (!i[1808]) | ( l_25 [3] &  i[1808]);
assign l_24[4]    = (!i[1808]) | ( l_25 [4] &  i[1808]);
assign l_24[5]    = ( l_25 [5] & !i[1808]);
assign l_24[6]    = ( l_25 [6] & !i[1808]);
assign l_24[7]    = (!i[1808]) | ( l_25 [7] &  i[1808]);
assign l_24[8]    = (!i[1808]) | ( l_25 [8] &  i[1808]);
assign l_24[9]    = ( l_25 [9] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[10]    = ( l_25 [10]);
assign l_24[11]    = ( l_25 [11] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[12]    = ( l_25 [10] & !i[1808]) | ( l_25 [12] &  i[1808]);
assign l_24[13]    = ( l_25 [10] & !i[1808]) | ( l_25 [13] &  i[1808]);
assign l_24[14]    = ( l_25 [14] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[15]    = ( l_25 [15] & !i[1808]) | ( l_25 [10] &  i[1808]);
assign l_24[16]    = ( l_25 [10] & !i[1808]) | ( l_25 [16] &  i[1808]);
assign l_24[17]    = ( l_25 [10] & !i[1808]) | ( l_25 [17] &  i[1808]);
assign l_24[18]    = ( l_25 [18]);
assign l_24[19]    = ( l_25 [19]);
assign l_24[20]    = ( l_25 [20]);
assign l_24[21]    = ( l_25 [21]);
assign l_24[22]    = ( l_25 [22]);
assign l_24[23]    = ( l_25 [23]);
assign l_24[24]    = ( l_25 [24]);
assign l_24[25]    = ( l_25 [25]);
assign l_24[26]    = ( l_25 [26]);
assign l_24[27]    = ( l_25 [27]);
assign l_24[28]    = ( l_25 [28]);
assign l_24[29]    = ( l_25 [29]);
assign l_24[30]    = ( l_25 [30]);
assign l_24[31]    = ( l_25 [31]);
assign l_24[32]    = ( l_25 [32]);
assign l_24[33]    = ( l_25 [33]);
assign l_24[34]    = ( l_25 [34]);
assign l_24[35]    = ( l_25 [35]);
assign l_24[36]    = ( l_25 [36]);
assign l_24[37]    = ( l_25 [37]);
assign l_24[38]    = ( l_25 [38]);
assign l_24[39]    = ( l_25 [39]);
assign l_24[40]    = ( l_25 [40]);
assign l_24[41]    = ( l_25 [41]);
assign l_24[42]    = ( l_25 [42]);
assign l_24[43]    = ( l_25 [43]);
assign l_24[44]    = ( l_25 [44]);
assign l_24[45]    = ( l_25 [45]);
assign l_24[46]    = ( l_25 [46]);
assign l_24[47]    = ( l_25 [47]);
assign l_24[48]    = ( l_25 [48]);
assign l_24[49]    = ( l_25 [49]);
assign l_24[50]    = ( l_25 [50] & !i[1808]) | ( l_25 [51] &  i[1808]);
assign l_24[51]    = ( l_25 [52] & !i[1808]) | ( l_25 [53] &  i[1808]);
assign l_25[0]    = ( l_26 [0]);
assign l_25[1]    = ( l_26 [1] & !i[1799]);
assign l_25[2]    = ( l_26 [2] & !i[1799]);
assign l_25[3]    = (!i[1799]) | ( l_26 [3] &  i[1799]);
assign l_25[4]    = (!i[1799]) | ( l_26 [4] &  i[1799]);
assign l_25[5]    = ( l_26 [5] & !i[1799]);
assign l_25[6]    = ( l_26 [6] & !i[1799]);
assign l_25[7]    = (!i[1799]) | ( l_26 [7] &  i[1799]);
assign l_25[8]    = (!i[1799]) | ( l_26 [8] &  i[1799]);
assign l_25[9]    = ( l_26 [9] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[10]    = ( l_26 [10]);
assign l_25[11]    = ( l_26 [11] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[12]    = ( l_26 [10] & !i[1799]) | ( l_26 [12] &  i[1799]);
assign l_25[13]    = ( l_26 [10] & !i[1799]) | ( l_26 [13] &  i[1799]);
assign l_25[14]    = ( l_26 [14] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[15]    = ( l_26 [15] & !i[1799]) | ( l_26 [10] &  i[1799]);
assign l_25[16]    = ( l_26 [10] & !i[1799]) | ( l_26 [16] &  i[1799]);
assign l_25[17]    = ( l_26 [10] & !i[1799]) | ( l_26 [17] &  i[1799]);
assign l_25[18]    = ( l_26 [18] & !i[1799]) | ( l_26 [19] &  i[1799]);
assign l_25[19]    = ( l_26 [20] & !i[1799]) | ( l_26 [21] &  i[1799]);
assign l_25[20]    = ( l_26 [22] & !i[1799]) | ( l_26 [23] &  i[1799]);
assign l_25[21]    = ( l_26 [24] & !i[1799]) | ( l_26 [25] &  i[1799]);
assign l_25[22]    = ( l_26 [26] & !i[1799]) | ( l_26 [27] &  i[1799]);
assign l_25[23]    = ( l_26 [28] & !i[1799]) | ( l_26 [29] &  i[1799]);
assign l_25[24]    = ( l_26 [30] & !i[1799]) | ( l_26 [31] &  i[1799]);
assign l_25[25]    = ( l_26 [32] & !i[1799]) | ( l_26 [33] &  i[1799]);
assign l_25[26]    = ( l_26 [34] & !i[1799]) | ( l_26 [35] &  i[1799]);
assign l_25[27]    = ( l_26 [36] & !i[1799]) | ( l_26 [37] &  i[1799]);
assign l_25[28]    = ( l_26 [38] & !i[1799]) | ( l_26 [39] &  i[1799]);
assign l_25[29]    = ( l_26 [40] & !i[1799]) | ( l_26 [41] &  i[1799]);
assign l_25[30]    = ( l_26 [42] & !i[1799]) | ( l_26 [43] &  i[1799]);
assign l_25[31]    = ( l_26 [44] & !i[1799]) | ( l_26 [45] &  i[1799]);
assign l_25[32]    = ( l_26 [46] & !i[1799]) | ( l_26 [47] &  i[1799]);
assign l_25[33]    = ( l_26 [48] & !i[1799]) | ( l_26 [49] &  i[1799]);
assign l_25[34]    = ( l_26 [50] & !i[1799]) | ( l_26 [51] &  i[1799]);
assign l_25[35]    = ( l_26 [52] & !i[1799]) | ( l_26 [53] &  i[1799]);
assign l_25[36]    = ( l_26 [54] & !i[1799]) | ( l_26 [55] &  i[1799]);
assign l_25[37]    = ( l_26 [56] & !i[1799]) | ( l_26 [57] &  i[1799]);
assign l_25[38]    = ( l_26 [58] & !i[1799]) | ( l_26 [59] &  i[1799]);
assign l_25[39]    = ( l_26 [60] & !i[1799]) | ( l_26 [61] &  i[1799]);
assign l_25[40]    = ( l_26 [62] & !i[1799]) | ( l_26 [63] &  i[1799]);
assign l_25[41]    = ( l_26 [64] & !i[1799]) | ( l_26 [65] &  i[1799]);
assign l_25[42]    = ( l_26 [66] & !i[1799]) | ( l_26 [67] &  i[1799]);
assign l_25[43]    = ( l_26 [68] & !i[1799]) | ( l_26 [69] &  i[1799]);
assign l_25[44]    = ( l_26 [70] & !i[1799]) | ( l_26 [71] &  i[1799]);
assign l_25[45]    = ( l_26 [72] & !i[1799]) | ( l_26 [73] &  i[1799]);
assign l_25[46]    = ( l_26 [74] & !i[1799]) | ( l_26 [75] &  i[1799]);
assign l_25[47]    = ( l_26 [76] & !i[1799]) | ( l_26 [77] &  i[1799]);
assign l_25[48]    = ( l_26 [78] & !i[1799]) | ( l_26 [79] &  i[1799]);
assign l_25[49]    = ( l_26 [80] & !i[1799]) | ( l_26 [81] &  i[1799]);
assign l_25[50]    = ( l_26 [82]);
assign l_25[51]    = ( l_26 [83]);
assign l_25[52]    = ( l_26 [84]);
assign l_25[53]    = ( l_26 [85]);
assign l_26[0]    = ( l_27 [0]);
assign l_26[1]    = ( l_27 [1] & !i[1802]);
assign l_26[2]    = ( l_27 [2] & !i[1802]);
assign l_26[3]    = (!i[1802]) | ( l_27 [3] &  i[1802]);
assign l_26[4]    = (!i[1802]) | ( l_27 [4] &  i[1802]);
assign l_26[5]    = ( l_27 [5] & !i[1802]);
assign l_26[6]    = ( l_27 [6] & !i[1802]);
assign l_26[7]    = (!i[1802]) | ( l_27 [7] &  i[1802]);
assign l_26[8]    = (!i[1802]) | ( l_27 [8] &  i[1802]);
assign l_26[9]    = ( l_27 [9] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[10]    = ( l_27 [10]);
assign l_26[11]    = ( l_27 [11] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[12]    = ( l_27 [10] & !i[1802]) | ( l_27 [12] &  i[1802]);
assign l_26[13]    = ( l_27 [10] & !i[1802]) | ( l_27 [13] &  i[1802]);
assign l_26[14]    = ( l_27 [14] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[15]    = ( l_27 [15] & !i[1802]) | ( l_27 [10] &  i[1802]);
assign l_26[16]    = ( l_27 [10] & !i[1802]) | ( l_27 [16] &  i[1802]);
assign l_26[17]    = ( l_27 [10] & !i[1802]) | ( l_27 [17] &  i[1802]);
assign l_26[18]    = ( l_27 [18]);
assign l_26[19]    = ( l_27 [19]);
assign l_26[20]    = ( l_27 [20]);
assign l_26[21]    = ( l_27 [21]);
assign l_26[22]    = ( l_27 [22]);
assign l_26[23]    = ( l_27 [23]);
assign l_26[24]    = ( l_27 [24]);
assign l_26[25]    = ( l_27 [25]);
assign l_26[26]    = ( l_27 [26]);
assign l_26[27]    = ( l_27 [27]);
assign l_26[28]    = ( l_27 [28]);
assign l_26[29]    = ( l_27 [29]);
assign l_26[30]    = ( l_27 [30]);
assign l_26[31]    = ( l_27 [31]);
assign l_26[32]    = ( l_27 [32]);
assign l_26[33]    = ( l_27 [33]);
assign l_26[34]    = ( l_27 [34]);
assign l_26[35]    = ( l_27 [35]);
assign l_26[36]    = ( l_27 [36]);
assign l_26[37]    = ( l_27 [37]);
assign l_26[38]    = ( l_27 [38]);
assign l_26[39]    = ( l_27 [39]);
assign l_26[40]    = ( l_27 [40]);
assign l_26[41]    = ( l_27 [41]);
assign l_26[42]    = ( l_27 [42]);
assign l_26[43]    = ( l_27 [43]);
assign l_26[44]    = ( l_27 [44]);
assign l_26[45]    = ( l_27 [45]);
assign l_26[46]    = ( l_27 [46]);
assign l_26[47]    = ( l_27 [47]);
assign l_26[48]    = ( l_27 [48]);
assign l_26[49]    = ( l_27 [49]);
assign l_26[50]    = ( l_27 [50]);
assign l_26[51]    = ( l_27 [51]);
assign l_26[52]    = ( l_27 [52]);
assign l_26[53]    = ( l_27 [53]);
assign l_26[54]    = ( l_27 [54]);
assign l_26[55]    = ( l_27 [55]);
assign l_26[56]    = ( l_27 [56]);
assign l_26[57]    = ( l_27 [57]);
assign l_26[58]    = ( l_27 [58]);
assign l_26[59]    = ( l_27 [59]);
assign l_26[60]    = ( l_27 [60]);
assign l_26[61]    = ( l_27 [61]);
assign l_26[62]    = ( l_27 [62]);
assign l_26[63]    = ( l_27 [63]);
assign l_26[64]    = ( l_27 [64]);
assign l_26[65]    = ( l_27 [65]);
assign l_26[66]    = ( l_27 [66]);
assign l_26[67]    = ( l_27 [67]);
assign l_26[68]    = ( l_27 [68]);
assign l_26[69]    = ( l_27 [69]);
assign l_26[70]    = ( l_27 [70]);
assign l_26[71]    = ( l_27 [71]);
assign l_26[72]    = ( l_27 [72]);
assign l_26[73]    = ( l_27 [73]);
assign l_26[74]    = ( l_27 [74]);
assign l_26[75]    = ( l_27 [75]);
assign l_26[76]    = ( l_27 [76]);
assign l_26[77]    = ( l_27 [77]);
assign l_26[78]    = ( l_27 [78]);
assign l_26[79]    = ( l_27 [79]);
assign l_26[80]    = ( l_27 [80]);
assign l_26[81]    = ( l_27 [81]);
assign l_26[82]    = ( l_27 [82] & !i[1802]) | ( l_27 [83] &  i[1802]);
assign l_26[83]    = ( l_27 [84] & !i[1802]) | ( l_27 [85] &  i[1802]);
assign l_26[84]    = ( l_27 [86] & !i[1802]) | ( l_27 [87] &  i[1802]);
assign l_26[85]    = ( l_27 [88] & !i[1802]) | ( l_27 [89] &  i[1802]);
assign l_27[0]    = ( l_28 [0]);
assign l_27[1]    = ( l_28 [1] & !i[1806]);
assign l_27[2]    = ( l_28 [2] & !i[1806]);
assign l_27[3]    = (!i[1806]) | ( l_28 [3] &  i[1806]);
assign l_27[4]    = (!i[1806]) | ( l_28 [4] &  i[1806]);
assign l_27[5]    = ( l_28 [5] & !i[1806]);
assign l_27[6]    = ( l_28 [6] & !i[1806]);
assign l_27[7]    = (!i[1806]) | ( l_28 [7] &  i[1806]);
assign l_27[8]    = (!i[1806]) | ( l_28 [8] &  i[1806]);
assign l_27[9]    = ( l_28 [9] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[10]    = ( l_28 [10]);
assign l_27[11]    = ( l_28 [11] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[12]    = ( l_28 [10] & !i[1806]) | ( l_28 [12] &  i[1806]);
assign l_27[13]    = ( l_28 [10] & !i[1806]) | ( l_28 [13] &  i[1806]);
assign l_27[14]    = ( l_28 [14] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[15]    = ( l_28 [15] & !i[1806]) | ( l_28 [10] &  i[1806]);
assign l_27[16]    = ( l_28 [10] & !i[1806]) | ( l_28 [16] &  i[1806]);
assign l_27[17]    = ( l_28 [10] & !i[1806]) | ( l_28 [17] &  i[1806]);
assign l_27[18]    = ( l_28 [18]);
assign l_27[19]    = ( l_28 [19]);
assign l_27[20]    = ( l_28 [20]);
assign l_27[21]    = ( l_28 [21]);
assign l_27[22]    = ( l_28 [22]);
assign l_27[23]    = ( l_28 [23]);
assign l_27[24]    = ( l_28 [24]);
assign l_27[25]    = ( l_28 [25]);
assign l_27[26]    = ( l_28 [26]);
assign l_27[27]    = ( l_28 [27]);
assign l_27[28]    = ( l_28 [28]);
assign l_27[29]    = ( l_28 [29]);
assign l_27[30]    = ( l_28 [30]);
assign l_27[31]    = ( l_28 [31]);
assign l_27[32]    = ( l_28 [32]);
assign l_27[33]    = ( l_28 [33]);
assign l_27[34]    = ( l_28 [34]);
assign l_27[35]    = ( l_28 [35]);
assign l_27[36]    = ( l_28 [36]);
assign l_27[37]    = ( l_28 [37]);
assign l_27[38]    = ( l_28 [38]);
assign l_27[39]    = ( l_28 [39]);
assign l_27[40]    = ( l_28 [40]);
assign l_27[41]    = ( l_28 [41]);
assign l_27[42]    = ( l_28 [42]);
assign l_27[43]    = ( l_28 [43]);
assign l_27[44]    = ( l_28 [44]);
assign l_27[45]    = ( l_28 [45]);
assign l_27[46]    = ( l_28 [46]);
assign l_27[47]    = ( l_28 [47]);
assign l_27[48]    = ( l_28 [48]);
assign l_27[49]    = ( l_28 [49]);
assign l_27[50]    = ( l_28 [50]);
assign l_27[51]    = ( l_28 [51]);
assign l_27[52]    = ( l_28 [52]);
assign l_27[53]    = ( l_28 [53]);
assign l_27[54]    = ( l_28 [54]);
assign l_27[55]    = ( l_28 [55]);
assign l_27[56]    = ( l_28 [56]);
assign l_27[57]    = ( l_28 [57]);
assign l_27[58]    = ( l_28 [58]);
assign l_27[59]    = ( l_28 [59]);
assign l_27[60]    = ( l_28 [60]);
assign l_27[61]    = ( l_28 [61]);
assign l_27[62]    = ( l_28 [62]);
assign l_27[63]    = ( l_28 [63]);
assign l_27[64]    = ( l_28 [64]);
assign l_27[65]    = ( l_28 [65]);
assign l_27[66]    = ( l_28 [66]);
assign l_27[67]    = ( l_28 [67]);
assign l_27[68]    = ( l_28 [68]);
assign l_27[69]    = ( l_28 [69]);
assign l_27[70]    = ( l_28 [70]);
assign l_27[71]    = ( l_28 [71]);
assign l_27[72]    = ( l_28 [72]);
assign l_27[73]    = ( l_28 [73]);
assign l_27[74]    = ( l_28 [74]);
assign l_27[75]    = ( l_28 [75]);
assign l_27[76]    = ( l_28 [76]);
assign l_27[77]    = ( l_28 [77]);
assign l_27[78]    = ( l_28 [78]);
assign l_27[79]    = ( l_28 [79]);
assign l_27[80]    = ( l_28 [80]);
assign l_27[81]    = ( l_28 [81]);
assign l_27[82]    = ( l_28 [82] & !i[1806]) | ( l_28 [83] &  i[1806]);
assign l_27[83]    = ( l_28 [84] & !i[1806]) | ( l_28 [85] &  i[1806]);
assign l_27[84]    = ( l_28 [86] & !i[1806]) | ( l_28 [87] &  i[1806]);
assign l_27[85]    = ( l_28 [88] & !i[1806]) | ( l_28 [89] &  i[1806]);
assign l_27[86]    = ( l_28 [90] & !i[1806]) | ( l_28 [91] &  i[1806]);
assign l_27[87]    = ( l_28 [92] & !i[1806]) | ( l_28 [93] &  i[1806]);
assign l_27[88]    = ( l_28 [94] & !i[1806]) | ( l_28 [95] &  i[1806]);
assign l_27[89]    = ( l_28 [96] & !i[1806]) | ( l_28 [97] &  i[1806]);
assign l_28[0]    = ( l_29 [0]);
assign l_28[1]    = ( l_29 [1] & !i[1816]);
assign l_28[2]    = ( l_29 [2] & !i[1816]);
assign l_28[3]    = (!i[1816]) | ( l_29 [3] &  i[1816]);
assign l_28[4]    = (!i[1816]) | ( l_29 [4] &  i[1816]);
assign l_28[5]    = ( l_29 [5] & !i[1816]);
assign l_28[6]    = ( l_29 [6] & !i[1816]);
assign l_28[7]    = (!i[1816]) | ( l_29 [7] &  i[1816]);
assign l_28[8]    = (!i[1816]) | ( l_29 [8] &  i[1816]);
assign l_28[9]    = ( l_29 [9] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[10]    = ( l_29 [10]);
assign l_28[11]    = ( l_29 [11] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[12]    = ( l_29 [10] & !i[1816]) | ( l_29 [12] &  i[1816]);
assign l_28[13]    = ( l_29 [10] & !i[1816]) | ( l_29 [13] &  i[1816]);
assign l_28[14]    = ( l_29 [14] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[15]    = ( l_29 [15] & !i[1816]) | ( l_29 [10] &  i[1816]);
assign l_28[16]    = ( l_29 [10] & !i[1816]) | ( l_29 [16] &  i[1816]);
assign l_28[17]    = ( l_29 [10] & !i[1816]) | ( l_29 [17] &  i[1816]);
assign l_28[18]    = ( l_29 [18]);
assign l_28[19]    = ( l_29 [19]);
assign l_28[20]    = ( l_29 [20]);
assign l_28[21]    = ( l_29 [21]);
assign l_28[22]    = ( l_29 [22]);
assign l_28[23]    = ( l_29 [23]);
assign l_28[24]    = ( l_29 [24]);
assign l_28[25]    = ( l_29 [25]);
assign l_28[26]    = ( l_29 [26]);
assign l_28[27]    = ( l_29 [27]);
assign l_28[28]    = ( l_29 [28]);
assign l_28[29]    = ( l_29 [29]);
assign l_28[30]    = ( l_29 [30]);
assign l_28[31]    = ( l_29 [31]);
assign l_28[32]    = ( l_29 [32]);
assign l_28[33]    = ( l_29 [33]);
assign l_28[34]    = ( l_29 [34]);
assign l_28[35]    = ( l_29 [35]);
assign l_28[36]    = ( l_29 [36]);
assign l_28[37]    = ( l_29 [37]);
assign l_28[38]    = ( l_29 [38]);
assign l_28[39]    = ( l_29 [39]);
assign l_28[40]    = ( l_29 [40]);
assign l_28[41]    = ( l_29 [41]);
assign l_28[42]    = ( l_29 [42]);
assign l_28[43]    = ( l_29 [43]);
assign l_28[44]    = ( l_29 [44]);
assign l_28[45]    = ( l_29 [45]);
assign l_28[46]    = ( l_29 [46]);
assign l_28[47]    = ( l_29 [47]);
assign l_28[48]    = ( l_29 [48]);
assign l_28[49]    = ( l_29 [49]);
assign l_28[50]    = ( l_29 [50]);
assign l_28[51]    = ( l_29 [51]);
assign l_28[52]    = ( l_29 [52]);
assign l_28[53]    = ( l_29 [53]);
assign l_28[54]    = ( l_29 [54]);
assign l_28[55]    = ( l_29 [55]);
assign l_28[56]    = ( l_29 [56]);
assign l_28[57]    = ( l_29 [57]);
assign l_28[58]    = ( l_29 [58]);
assign l_28[59]    = ( l_29 [59]);
assign l_28[60]    = ( l_29 [60]);
assign l_28[61]    = ( l_29 [61]);
assign l_28[62]    = ( l_29 [62]);
assign l_28[63]    = ( l_29 [63]);
assign l_28[64]    = ( l_29 [64]);
assign l_28[65]    = ( l_29 [65]);
assign l_28[66]    = ( l_29 [66]);
assign l_28[67]    = ( l_29 [67]);
assign l_28[68]    = ( l_29 [68]);
assign l_28[69]    = ( l_29 [69]);
assign l_28[70]    = ( l_29 [70]);
assign l_28[71]    = ( l_29 [71]);
assign l_28[72]    = ( l_29 [72]);
assign l_28[73]    = ( l_29 [73]);
assign l_28[74]    = ( l_29 [74]);
assign l_28[75]    = ( l_29 [75]);
assign l_28[76]    = ( l_29 [76]);
assign l_28[77]    = ( l_29 [77]);
assign l_28[78]    = ( l_29 [78]);
assign l_28[79]    = ( l_29 [79]);
assign l_28[80]    = ( l_29 [80]);
assign l_28[81]    = ( l_29 [81]);
assign l_28[82]    = ( l_29 [82] & !i[1816]) | ( l_29 [83] &  i[1816]);
assign l_28[83]    = ( l_29 [84] & !i[1816]) | ( l_29 [85] &  i[1816]);
assign l_28[84]    = ( l_29 [86] & !i[1816]) | ( l_29 [87] &  i[1816]);
assign l_28[85]    = ( l_29 [88] & !i[1816]) | ( l_29 [89] &  i[1816]);
assign l_28[86]    = ( l_29 [90] & !i[1816]) | ( l_29 [91] &  i[1816]);
assign l_28[87]    = ( l_29 [92] & !i[1816]) | ( l_29 [93] &  i[1816]);
assign l_28[88]    = ( l_29 [94] & !i[1816]) | ( l_29 [95] &  i[1816]);
assign l_28[89]    = ( l_29 [96] & !i[1816]) | ( l_29 [97] &  i[1816]);
assign l_28[90]    = ( l_29 [98] & !i[1816]) | ( l_29 [99] &  i[1816]);
assign l_28[91]    = ( l_29 [100] & !i[1816]) | ( l_29 [101] &  i[1816]);
assign l_28[92]    = ( l_29 [102] & !i[1816]) | ( l_29 [103] &  i[1816]);
assign l_28[93]    = ( l_29 [104] & !i[1816]) | ( l_29 [105] &  i[1816]);
assign l_28[94]    = ( l_29 [106] & !i[1816]) | ( l_29 [107] &  i[1816]);
assign l_28[95]    = ( l_29 [108] & !i[1816]) | ( l_29 [109] &  i[1816]);
assign l_28[96]    = ( l_29 [110] & !i[1816]) | ( l_29 [111] &  i[1816]);
assign l_28[97]    = ( l_29 [112] & !i[1816]) | ( l_29 [113] &  i[1816]);
assign l_29[0]    = ( l_30 [0]);
assign l_29[1]    = ( l_30 [1] & !i[1810]);
assign l_29[2]    = ( l_30 [2] & !i[1810]);
assign l_29[3]    = (!i[1810]) | ( l_30 [3] &  i[1810]);
assign l_29[4]    = (!i[1810]) | ( l_30 [4] &  i[1810]);
assign l_29[5]    = ( l_30 [5] & !i[1810]);
assign l_29[6]    = ( l_30 [6] & !i[1810]);
assign l_29[7]    = (!i[1810]) | ( l_30 [7] &  i[1810]);
assign l_29[8]    = (!i[1810]) | ( l_30 [8] &  i[1810]);
assign l_29[9]    = ( l_30 [9] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[10]    = ( l_30 [10]);
assign l_29[11]    = ( l_30 [11] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[12]    = ( l_30 [10] & !i[1810]) | ( l_30 [12] &  i[1810]);
assign l_29[13]    = ( l_30 [10] & !i[1810]) | ( l_30 [13] &  i[1810]);
assign l_29[14]    = ( l_30 [14] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[15]    = ( l_30 [15] & !i[1810]) | ( l_30 [10] &  i[1810]);
assign l_29[16]    = ( l_30 [10] & !i[1810]) | ( l_30 [16] &  i[1810]);
assign l_29[17]    = ( l_30 [10] & !i[1810]) | ( l_30 [17] &  i[1810]);
assign l_29[18]    = ( l_30 [18]);
assign l_29[19]    = ( l_30 [19]);
assign l_29[20]    = ( l_30 [20]);
assign l_29[21]    = ( l_30 [21]);
assign l_29[22]    = ( l_30 [22]);
assign l_29[23]    = ( l_30 [23]);
assign l_29[24]    = ( l_30 [24]);
assign l_29[25]    = ( l_30 [25]);
assign l_29[26]    = ( l_30 [26]);
assign l_29[27]    = ( l_30 [27]);
assign l_29[28]    = ( l_30 [28]);
assign l_29[29]    = ( l_30 [29]);
assign l_29[30]    = ( l_30 [30]);
assign l_29[31]    = ( l_30 [31]);
assign l_29[32]    = ( l_30 [32]);
assign l_29[33]    = ( l_30 [33]);
assign l_29[34]    = ( l_30 [34]);
assign l_29[35]    = ( l_30 [35]);
assign l_29[36]    = ( l_30 [36]);
assign l_29[37]    = ( l_30 [37]);
assign l_29[38]    = ( l_30 [38]);
assign l_29[39]    = ( l_30 [39]);
assign l_29[40]    = ( l_30 [40]);
assign l_29[41]    = ( l_30 [41]);
assign l_29[42]    = ( l_30 [42]);
assign l_29[43]    = ( l_30 [43]);
assign l_29[44]    = ( l_30 [44]);
assign l_29[45]    = ( l_30 [45]);
assign l_29[46]    = ( l_30 [46]);
assign l_29[47]    = ( l_30 [47]);
assign l_29[48]    = ( l_30 [48]);
assign l_29[49]    = ( l_30 [49]);
assign l_29[50]    = ( l_30 [50]);
assign l_29[51]    = ( l_30 [51]);
assign l_29[52]    = ( l_30 [52]);
assign l_29[53]    = ( l_30 [53]);
assign l_29[54]    = ( l_30 [54]);
assign l_29[55]    = ( l_30 [55]);
assign l_29[56]    = ( l_30 [56]);
assign l_29[57]    = ( l_30 [57]);
assign l_29[58]    = ( l_30 [58]);
assign l_29[59]    = ( l_30 [59]);
assign l_29[60]    = ( l_30 [60]);
assign l_29[61]    = ( l_30 [61]);
assign l_29[62]    = ( l_30 [62]);
assign l_29[63]    = ( l_30 [63]);
assign l_29[64]    = ( l_30 [64]);
assign l_29[65]    = ( l_30 [65]);
assign l_29[66]    = ( l_30 [66]);
assign l_29[67]    = ( l_30 [67]);
assign l_29[68]    = ( l_30 [68]);
assign l_29[69]    = ( l_30 [69]);
assign l_29[70]    = ( l_30 [70]);
assign l_29[71]    = ( l_30 [71]);
assign l_29[72]    = ( l_30 [72]);
assign l_29[73]    = ( l_30 [73]);
assign l_29[74]    = ( l_30 [74]);
assign l_29[75]    = ( l_30 [75]);
assign l_29[76]    = ( l_30 [76]);
assign l_29[77]    = ( l_30 [77]);
assign l_29[78]    = ( l_30 [78]);
assign l_29[79]    = ( l_30 [79]);
assign l_29[80]    = ( l_30 [80]);
assign l_29[81]    = ( l_30 [81]);
assign l_29[82]    = ( l_30 [82] & !i[1810]) | ( l_30 [83] &  i[1810]);
assign l_29[83]    = ( l_30 [84] & !i[1810]) | ( l_30 [85] &  i[1810]);
assign l_29[84]    = ( l_30 [86] & !i[1810]) | ( l_30 [87] &  i[1810]);
assign l_29[85]    = ( l_30 [88] & !i[1810]) | ( l_30 [89] &  i[1810]);
assign l_29[86]    = ( l_30 [90] & !i[1810]) | ( l_30 [91] &  i[1810]);
assign l_29[87]    = ( l_30 [92] & !i[1810]) | ( l_30 [93] &  i[1810]);
assign l_29[88]    = ( l_30 [94] & !i[1810]) | ( l_30 [95] &  i[1810]);
assign l_29[89]    = ( l_30 [96] & !i[1810]) | ( l_30 [97] &  i[1810]);
assign l_29[90]    = ( l_30 [98] & !i[1810]) | ( l_30 [99] &  i[1810]);
assign l_29[91]    = ( l_30 [100] & !i[1810]) | ( l_30 [101] &  i[1810]);
assign l_29[92]    = ( l_30 [102] & !i[1810]) | ( l_30 [103] &  i[1810]);
assign l_29[93]    = ( l_30 [104] & !i[1810]) | ( l_30 [105] &  i[1810]);
assign l_29[94]    = ( l_30 [106] & !i[1810]) | ( l_30 [107] &  i[1810]);
assign l_29[95]    = ( l_30 [108] & !i[1810]) | ( l_30 [109] &  i[1810]);
assign l_29[96]    = ( l_30 [110] & !i[1810]) | ( l_30 [111] &  i[1810]);
assign l_29[97]    = ( l_30 [112] & !i[1810]) | ( l_30 [113] &  i[1810]);
assign l_29[98]    = ( l_30 [114] & !i[1810]) | ( l_30 [115] &  i[1810]);
assign l_29[99]    = ( l_30 [116] & !i[1810]) | ( l_30 [117] &  i[1810]);
assign l_29[100]    = ( l_30 [118] & !i[1810]) | ( l_30 [119] &  i[1810]);
assign l_29[101]    = ( l_30 [120] & !i[1810]) | ( l_30 [121] &  i[1810]);
assign l_29[102]    = ( l_30 [122] & !i[1810]) | ( l_30 [123] &  i[1810]);
assign l_29[103]    = ( l_30 [124] & !i[1810]) | ( l_30 [125] &  i[1810]);
assign l_29[104]    = ( l_30 [126] & !i[1810]) | ( l_30 [127] &  i[1810]);
assign l_29[105]    = ( l_30 [128] & !i[1810]) | ( l_30 [129] &  i[1810]);
assign l_29[106]    = ( l_30 [130] & !i[1810]) | ( l_30 [131] &  i[1810]);
assign l_29[107]    = ( l_30 [132] & !i[1810]) | ( l_30 [133] &  i[1810]);
assign l_29[108]    = ( l_30 [134] & !i[1810]) | ( l_30 [135] &  i[1810]);
assign l_29[109]    = ( l_30 [136] & !i[1810]) | ( l_30 [137] &  i[1810]);
assign l_29[110]    = ( l_30 [138] & !i[1810]) | ( l_30 [139] &  i[1810]);
assign l_29[111]    = ( l_30 [140] & !i[1810]) | ( l_30 [141] &  i[1810]);
assign l_29[112]    = ( l_30 [142] & !i[1810]) | ( l_30 [143] &  i[1810]);
assign l_29[113]    = ( l_30 [144] & !i[1810]) | ( l_30 [145] &  i[1810]);

endmodule
